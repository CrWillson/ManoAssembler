
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.0 | 2017-01-18 18:54:33</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-103.148,1.08472,199.294,-151.665</PageViewport>
<gate>
<ID>2</ID>
<type>AM_REGISTER16</type>
<position>25.5,-78.5</position>
<input>
<ID>IN_0</ID>214 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_10</ID>221 </input>
<input>
<ID>IN_11</ID>225 </input>
<input>
<ID>IN_12</ID>222 </input>
<input>
<ID>IN_13</ID>217 </input>
<input>
<ID>IN_14</ID>218 </input>
<input>
<ID>IN_15</ID>210 </input>
<input>
<ID>IN_2</ID>223 </input>
<input>
<ID>IN_3</ID>220 </input>
<input>
<ID>IN_4</ID>213 </input>
<input>
<ID>IN_5</ID>215 </input>
<input>
<ID>IN_6</ID>224 </input>
<input>
<ID>IN_7</ID>211 </input>
<input>
<ID>IN_8</ID>212 </input>
<input>
<ID>IN_9</ID>216 </input>
<output>
<ID>OUT_0</ID>547 </output>
<output>
<ID>OUT_1</ID>548 </output>
<output>
<ID>OUT_10</ID>557 </output>
<output>
<ID>OUT_11</ID>558 </output>
<output>
<ID>OUT_12</ID>559 </output>
<output>
<ID>OUT_13</ID>560 </output>
<output>
<ID>OUT_14</ID>561 </output>
<output>
<ID>OUT_15</ID>562 </output>
<output>
<ID>OUT_2</ID>549 </output>
<output>
<ID>OUT_3</ID>550 </output>
<output>
<ID>OUT_4</ID>551 </output>
<output>
<ID>OUT_5</ID>552 </output>
<output>
<ID>OUT_6</ID>553 </output>
<output>
<ID>OUT_7</ID>554 </output>
<output>
<ID>OUT_8</ID>555 </output>
<output>
<ID>OUT_9</ID>556 </output>
<input>
<ID>clear</ID>582 </input>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>count_enable</ID>581 </input>
<input>
<ID>load</ID>580 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>10</ID>
<type>AI_REGISTER12</type>
<position>25.5,-46.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_10</ID>39 </input>
<input>
<ID>IN_11</ID>40 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>30 </input>
<input>
<ID>IN_4</ID>33 </input>
<input>
<ID>IN_5</ID>34 </input>
<input>
<ID>IN_6</ID>35 </input>
<input>
<ID>IN_7</ID>36 </input>
<input>
<ID>IN_8</ID>37 </input>
<input>
<ID>IN_9</ID>38 </input>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>12 </output>
<output>
<ID>OUT_10</ID>3 </output>
<output>
<ID>OUT_11</ID>2 </output>
<output>
<ID>OUT_2</ID>11 </output>
<output>
<ID>OUT_3</ID>10 </output>
<output>
<ID>OUT_4</ID>9 </output>
<output>
<ID>OUT_5</ID>8 </output>
<output>
<ID>OUT_6</ID>7 </output>
<output>
<ID>OUT_7</ID>6 </output>
<output>
<ID>OUT_8</ID>5 </output>
<output>
<ID>OUT_9</ID>4 </output>
<input>
<ID>clear</ID>544 </input>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>count_enable</ID>543 </input>
<input>
<ID>load</ID>542 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>18</ID>
<type>BX_16X1_BUS_END</type>
<position>67,-44.5</position>
<input>
<ID>Bus_in_0</ID>41 </input>
<input>
<ID>IN_1</ID>42 </input>
<input>
<ID>IN_10</ID>56 </input>
<input>
<ID>IN_11</ID>50 </input>
<input>
<ID>IN_12</ID>51 </input>
<input>
<ID>IN_13</ID>54 </input>
<input>
<ID>IN_14</ID>55 </input>
<input>
<ID>IN_15</ID>53 </input>
<input>
<ID>IN_2</ID>47 </input>
<input>
<ID>IN_3</ID>43 </input>
<input>
<ID>IN_4</ID>44 </input>
<input>
<ID>IN_5</ID>45 </input>
<input>
<ID>IN_6</ID>48 </input>
<input>
<ID>IN_7</ID>46 </input>
<input>
<ID>IN_8</ID>49 </input>
<input>
<ID>IN_9</ID>52 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>8</ID>
<type>AI_RAM_12x16</type>
<position>74,-12</position>
<input>
<ID>ADDRESS_0</ID>1 </input>
<input>
<ID>ADDRESS_1</ID>12 </input>
<input>
<ID>ADDRESS_10</ID>3 </input>
<input>
<ID>ADDRESS_11</ID>2 </input>
<input>
<ID>ADDRESS_2</ID>11 </input>
<input>
<ID>ADDRESS_3</ID>10 </input>
<input>
<ID>ADDRESS_4</ID>9 </input>
<input>
<ID>ADDRESS_5</ID>8 </input>
<input>
<ID>ADDRESS_6</ID>7 </input>
<input>
<ID>ADDRESS_7</ID>6 </input>
<input>
<ID>ADDRESS_8</ID>5 </input>
<input>
<ID>ADDRESS_9</ID>4 </input>
<input>
<ID>DATA_IN_0</ID>58 </input>
<input>
<ID>DATA_IN_1</ID>59 </input>
<input>
<ID>DATA_IN_10</ID>68 </input>
<input>
<ID>DATA_IN_11</ID>69 </input>
<input>
<ID>DATA_IN_12</ID>60 </input>
<input>
<ID>DATA_IN_13</ID>62 </input>
<input>
<ID>DATA_IN_14</ID>72 </input>
<input>
<ID>DATA_IN_15</ID>70 </input>
<input>
<ID>DATA_IN_2</ID>57 </input>
<input>
<ID>DATA_IN_3</ID>63 </input>
<input>
<ID>DATA_IN_4</ID>64 </input>
<input>
<ID>DATA_IN_5</ID>61 </input>
<input>
<ID>DATA_IN_6</ID>65 </input>
<input>
<ID>DATA_IN_7</ID>66 </input>
<input>
<ID>DATA_IN_8</ID>71 </input>
<input>
<ID>DATA_IN_9</ID>67 </input>
<output>
<ID>DATA_OUT_0</ID>58 </output>
<output>
<ID>DATA_OUT_1</ID>59 </output>
<output>
<ID>DATA_OUT_10</ID>68 </output>
<output>
<ID>DATA_OUT_11</ID>69 </output>
<output>
<ID>DATA_OUT_12</ID>60 </output>
<output>
<ID>DATA_OUT_13</ID>62 </output>
<output>
<ID>DATA_OUT_14</ID>72 </output>
<output>
<ID>DATA_OUT_15</ID>70 </output>
<output>
<ID>DATA_OUT_2</ID>57 </output>
<output>
<ID>DATA_OUT_3</ID>63 </output>
<output>
<ID>DATA_OUT_4</ID>64 </output>
<output>
<ID>DATA_OUT_5</ID>61 </output>
<output>
<ID>DATA_OUT_6</ID>65 </output>
<output>
<ID>DATA_OUT_7</ID>66 </output>
<output>
<ID>DATA_OUT_8</ID>71 </output>
<output>
<ID>DATA_OUT_9</ID>67 </output>
<input>
<ID>ENABLE_0</ID>708 </input>
<input>
<ID>write_clock</ID>513 </input>
<input>
<ID>write_enable</ID>662 </input>
<gparam>angle 0.0</gparam>
<lparam>ADDRESS_BITS 12</lparam>
<lparam>DATA_BITS 16</lparam>
<lparam>Address:0 16640</lparam>
<lparam>Address:256 8459</lparam>
<lparam>Address:257 12556</lparam>
<lparam>Address:258 8461</lparam>
<lparam>Address:259 12558</lparam>
<lparam>Address:260 30720</lparam>
<lparam>Address:261 37132</lparam>
<lparam>Address:262 24844</lparam>
<lparam>Address:263 24846</lparam>
<lparam>Address:264 16645</lparam>
<lparam>Address:265 12559</lparam>
<lparam>Address:266 28673</lparam>
<lparam>Address:267 336</lparam>
<lparam>Address:268 346</lparam>
<lparam>Address:269 65526</lparam>
<lparam>Address:271 575</lparam>
<lparam>Address:336 25</lparam>
<lparam>Address:337 50</lparam>
<lparam>Address:338 75</lparam>
<lparam>Address:339 100</lparam>
<lparam>Address:340 25</lparam>
<lparam>Address:341 50</lparam>
<lparam>Address:342 75</lparam>
<lparam>Address:343 100</lparam>
<lparam>Address:344 25</lparam>
<lparam>Address:345 50</lparam></gate>
<gate>
<ID>16</ID>
<type>BX_16X1_BUS_END</type>
<position>17.5,-44.5</position>
<input>
<ID>Bus_in_0</ID>31 </input>
<input>
<ID>IN_1</ID>29 </input>
<input>
<ID>IN_10</ID>39 </input>
<input>
<ID>IN_11</ID>40 </input>
<input>
<ID>IN_2</ID>32 </input>
<input>
<ID>IN_3</ID>30 </input>
<input>
<ID>IN_4</ID>33 </input>
<input>
<ID>IN_5</ID>34 </input>
<input>
<ID>IN_6</ID>35 </input>
<input>
<ID>IN_7</ID>36 </input>
<input>
<ID>IN_8</ID>37 </input>
<input>
<ID>IN_9</ID>38 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>20</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>56,-44.5</position>
<input>
<ID>ENABLE_0</ID>545 </input>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>12 </input>
<input>
<ID>IN_10</ID>3 </input>
<input>
<ID>IN_11</ID>2 </input>
<input>
<ID>IN_2</ID>11 </input>
<input>
<ID>IN_3</ID>10 </input>
<input>
<ID>IN_4</ID>9 </input>
<input>
<ID>IN_5</ID>8 </input>
<input>
<ID>IN_6</ID>7 </input>
<input>
<ID>IN_7</ID>6 </input>
<input>
<ID>IN_8</ID>5 </input>
<input>
<ID>IN_9</ID>4 </input>
<output>
<ID>OUT_0</ID>41 </output>
<output>
<ID>OUT_1</ID>42 </output>
<output>
<ID>OUT_10</ID>56 </output>
<output>
<ID>OUT_11</ID>50 </output>
<output>
<ID>OUT_12</ID>51 </output>
<output>
<ID>OUT_13</ID>54 </output>
<output>
<ID>OUT_14</ID>55 </output>
<output>
<ID>OUT_15</ID>53 </output>
<output>
<ID>OUT_2</ID>47 </output>
<output>
<ID>OUT_3</ID>43 </output>
<output>
<ID>OUT_4</ID>44 </output>
<output>
<ID>OUT_5</ID>45 </output>
<output>
<ID>OUT_6</ID>48 </output>
<output>
<ID>OUT_7</ID>46 </output>
<output>
<ID>OUT_8</ID>49 </output>
<output>
<ID>OUT_9</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>22</ID>
<type>BX_16X1_BUS_END</type>
<position>81,-44.5</position>
<input>
<ID>Bus_in_0</ID>307 </input>
<input>
<ID>IN_1</ID>308 </input>
<input>
<ID>IN_10</ID>316 </input>
<input>
<ID>IN_11</ID>317 </input>
<input>
<ID>IN_2</ID>306 </input>
<input>
<ID>IN_3</ID>309 </input>
<input>
<ID>IN_4</ID>310 </input>
<input>
<ID>IN_5</ID>311 </input>
<input>
<ID>IN_6</ID>312 </input>
<input>
<ID>IN_7</ID>313 </input>
<input>
<ID>IN_8</ID>314 </input>
<input>
<ID>IN_9</ID>315 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>29</ID>
<type>AM_REGISTER16</type>
<position>25.5,-119.5</position>
<input>
<ID>IN_0</ID>237 </input>
<input>
<ID>IN_1</ID>226 </input>
<input>
<ID>IN_10</ID>240 </input>
<input>
<ID>IN_11</ID>228 </input>
<input>
<ID>IN_12</ID>229 </input>
<input>
<ID>IN_13</ID>241 </input>
<input>
<ID>IN_14</ID>234 </input>
<input>
<ID>IN_15</ID>230 </input>
<input>
<ID>IN_2</ID>236 </input>
<input>
<ID>IN_3</ID>227 </input>
<input>
<ID>IN_4</ID>235 </input>
<input>
<ID>IN_5</ID>238 </input>
<input>
<ID>IN_6</ID>232 </input>
<input>
<ID>IN_7</ID>239 </input>
<input>
<ID>IN_8</ID>231 </input>
<input>
<ID>IN_9</ID>233 </input>
<output>
<ID>OUT_0</ID>285 </output>
<output>
<ID>OUT_1</ID>274 </output>
<output>
<ID>OUT_10</ID>283 </output>
<output>
<ID>OUT_11</ID>284 </output>
<output>
<ID>OUT_12</ID>286 </output>
<output>
<ID>OUT_13</ID>288 </output>
<output>
<ID>OUT_14</ID>287 </output>
<output>
<ID>OUT_15</ID>289 </output>
<output>
<ID>OUT_2</ID>275 </output>
<output>
<ID>OUT_3</ID>276 </output>
<output>
<ID>OUT_4</ID>277 </output>
<output>
<ID>OUT_5</ID>278 </output>
<output>
<ID>OUT_6</ID>279 </output>
<output>
<ID>OUT_7</ID>280 </output>
<output>
<ID>OUT_8</ID>281 </output>
<output>
<ID>OUT_9</ID>282 </output>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>load</ID>584 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>223</ID>
<type>DA_FROM</type>
<position>52.5,-68</position>
<input>
<ID>IN_0</ID>583 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_bus</lparam></gate>
<gate>
<ID>31</ID>
<type>BX_16X1_BUS_END</type>
<position>67,-78.5</position>
<input>
<ID>Bus_in_0</ID>114 </input>
<input>
<ID>IN_1</ID>115 </input>
<input>
<ID>IN_10</ID>129 </input>
<input>
<ID>IN_11</ID>123 </input>
<input>
<ID>IN_12</ID>124 </input>
<input>
<ID>IN_13</ID>127 </input>
<input>
<ID>IN_14</ID>128 </input>
<input>
<ID>IN_15</ID>126 </input>
<input>
<ID>IN_2</ID>120 </input>
<input>
<ID>IN_3</ID>116 </input>
<input>
<ID>IN_4</ID>117 </input>
<input>
<ID>IN_5</ID>118 </input>
<input>
<ID>IN_6</ID>121 </input>
<input>
<ID>IN_7</ID>119 </input>
<input>
<ID>IN_8</ID>122 </input>
<input>
<ID>IN_9</ID>125 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>32</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>56,-78.5</position>
<input>
<ID>ENABLE_0</ID>583 </input>
<input>
<ID>IN_0</ID>547 </input>
<input>
<ID>IN_1</ID>548 </input>
<input>
<ID>IN_10</ID>557 </input>
<input>
<ID>IN_11</ID>558 </input>
<input>
<ID>IN_12</ID>559 </input>
<input>
<ID>IN_13</ID>560 </input>
<input>
<ID>IN_14</ID>561 </input>
<input>
<ID>IN_15</ID>562 </input>
<input>
<ID>IN_2</ID>549 </input>
<input>
<ID>IN_3</ID>550 </input>
<input>
<ID>IN_4</ID>551 </input>
<input>
<ID>IN_5</ID>552 </input>
<input>
<ID>IN_6</ID>553 </input>
<input>
<ID>IN_7</ID>554 </input>
<input>
<ID>IN_8</ID>555 </input>
<input>
<ID>IN_9</ID>556 </input>
<output>
<ID>OUT_0</ID>114 </output>
<output>
<ID>OUT_1</ID>115 </output>
<output>
<ID>OUT_10</ID>129 </output>
<output>
<ID>OUT_11</ID>123 </output>
<output>
<ID>OUT_12</ID>124 </output>
<output>
<ID>OUT_13</ID>127 </output>
<output>
<ID>OUT_14</ID>128 </output>
<output>
<ID>OUT_15</ID>126 </output>
<output>
<ID>OUT_2</ID>120 </output>
<output>
<ID>OUT_3</ID>116 </output>
<output>
<ID>OUT_4</ID>117 </output>
<output>
<ID>OUT_5</ID>118 </output>
<output>
<ID>OUT_6</ID>121 </output>
<output>
<ID>OUT_7</ID>119 </output>
<output>
<ID>OUT_8</ID>122 </output>
<output>
<ID>OUT_9</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>225</ID>
<type>DA_FROM</type>
<position>22.5,-108.5</position>
<input>
<ID>IN_0</ID>584 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR_LD</lparam></gate>
<gate>
<ID>97</ID>
<type>BB_CLOCK</type>
<position>-56.5,-60.5</position>
<output>
<ID>CLK</ID>486 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 3</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>86,-108.5</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_LD</lparam></gate>
<gate>
<ID>35</ID>
<type>BX_16X1_BUS_END</type>
<position>67,-119.5</position>
<input>
<ID>Bus_in_0</ID>162 </input>
<input>
<ID>IN_1</ID>163 </input>
<input>
<ID>IN_10</ID>177 </input>
<input>
<ID>IN_11</ID>171 </input>
<input>
<ID>IN_12</ID>172 </input>
<input>
<ID>IN_13</ID>175 </input>
<input>
<ID>IN_14</ID>176 </input>
<input>
<ID>IN_15</ID>174 </input>
<input>
<ID>IN_2</ID>168 </input>
<input>
<ID>IN_3</ID>164 </input>
<input>
<ID>IN_4</ID>165 </input>
<input>
<ID>IN_5</ID>166 </input>
<input>
<ID>IN_6</ID>169 </input>
<input>
<ID>IN_7</ID>167 </input>
<input>
<ID>IN_8</ID>170 </input>
<input>
<ID>IN_9</ID>173 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>99</ID>
<type>CC_PULSE</type>
<position>-56.5,-65.5</position>
<output>
<ID>OUT_0</ID>487 </output>
<gparam>CLICK_BOX -0.75,-0.75,0.75,0.75</gparam>
<gparam>PULSE_WIDTH 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>DA_FROM</type>
<position>22.5,-34.5</position>
<input>
<ID>IN_0</ID>542 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_LD</lparam></gate>
<gate>
<ID>36</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>56,-119.5</position>
<input>
<ID>ENABLE_0</ID>192 </input>
<input>
<ID>IN_0</ID>285 </input>
<input>
<ID>IN_1</ID>274 </input>
<input>
<ID>IN_10</ID>283 </input>
<input>
<ID>IN_11</ID>284 </input>
<input>
<ID>IN_12</ID>286 </input>
<input>
<ID>IN_13</ID>288 </input>
<input>
<ID>IN_14</ID>287 </input>
<input>
<ID>IN_15</ID>289 </input>
<input>
<ID>IN_2</ID>275 </input>
<input>
<ID>IN_3</ID>276 </input>
<input>
<ID>IN_4</ID>277 </input>
<input>
<ID>IN_5</ID>278 </input>
<input>
<ID>IN_6</ID>279 </input>
<input>
<ID>IN_7</ID>280 </input>
<input>
<ID>IN_8</ID>281 </input>
<input>
<ID>IN_9</ID>282 </input>
<output>
<ID>OUT_0</ID>162 </output>
<output>
<ID>OUT_1</ID>163 </output>
<output>
<ID>OUT_10</ID>177 </output>
<output>
<ID>OUT_11</ID>171 </output>
<output>
<ID>OUT_12</ID>172 </output>
<output>
<ID>OUT_13</ID>175 </output>
<output>
<ID>OUT_14</ID>176 </output>
<output>
<ID>OUT_15</ID>174 </output>
<output>
<ID>OUT_2</ID>168 </output>
<output>
<ID>OUT_3</ID>164 </output>
<output>
<ID>OUT_4</ID>165 </output>
<output>
<ID>OUT_5</ID>166 </output>
<output>
<ID>OUT_6</ID>169 </output>
<output>
<ID>OUT_7</ID>167 </output>
<output>
<ID>OUT_8</ID>170 </output>
<output>
<ID>OUT_9</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1097</ID>
<type>DE_TO</type>
<position>-41,-99</position>
<input>
<ID>IN_0</ID>1221 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR7</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>86,-106</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_INC</lparam></gate>
<gate>
<ID>101</ID>
<type>AA_MUX_2x1</type>
<position>-49,-63</position>
<input>
<ID>IN_0</ID>487 </input>
<input>
<ID>IN_1</ID>486 </input>
<output>
<ID>OUT</ID>489 </output>
<input>
<ID>SEL_0</ID>488 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>165</ID>
<type>DA_FROM</type>
<position>22.5,-32</position>
<input>
<ID>IN_0</ID>543 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_INC</lparam></gate>
<gate>
<ID>1092</ID>
<type>DE_TO</type>
<position>-50,-102</position>
<input>
<ID>IN_0</ID>1216 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR4</lparam></gate>
<gate>
<ID>40</ID>
<type>BX_16X1_BUS_END</type>
<position>17.5,-78.5</position>
<input>
<ID>Bus_in_0</ID>214 </input>
<input>
<ID>IN_1</ID>219 </input>
<input>
<ID>IN_10</ID>221 </input>
<input>
<ID>IN_11</ID>225 </input>
<input>
<ID>IN_12</ID>222 </input>
<input>
<ID>IN_13</ID>217 </input>
<input>
<ID>IN_14</ID>218 </input>
<input>
<ID>IN_15</ID>210 </input>
<input>
<ID>IN_2</ID>223 </input>
<input>
<ID>IN_3</ID>220 </input>
<input>
<ID>IN_4</ID>213 </input>
<input>
<ID>IN_5</ID>215 </input>
<input>
<ID>IN_6</ID>224 </input>
<input>
<ID>IN_7</ID>211 </input>
<input>
<ID>IN_8</ID>212 </input>
<input>
<ID>IN_9</ID>216 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>1093</ID>
<type>DE_TO</type>
<position>-41,-105</position>
<input>
<ID>IN_0</ID>1219 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR1</lparam></gate>
<gate>
<ID>41</ID>
<type>BX_16X1_BUS_END</type>
<position>17.5,-119.5</position>
<input>
<ID>Bus_in_0</ID>237 </input>
<input>
<ID>IN_1</ID>226 </input>
<input>
<ID>IN_10</ID>240 </input>
<input>
<ID>IN_11</ID>228 </input>
<input>
<ID>IN_12</ID>229 </input>
<input>
<ID>IN_13</ID>241 </input>
<input>
<ID>IN_14</ID>234 </input>
<input>
<ID>IN_15</ID>230 </input>
<input>
<ID>IN_2</ID>236 </input>
<input>
<ID>IN_3</ID>227 </input>
<input>
<ID>IN_4</ID>235 </input>
<input>
<ID>IN_5</ID>238 </input>
<input>
<ID>IN_6</ID>232 </input>
<input>
<ID>IN_7</ID>239 </input>
<input>
<ID>IN_8</ID>231 </input>
<input>
<ID>IN_9</ID>233 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>-44,-63</position>
<input>
<ID>IN_0</ID>489 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>169</ID>
<type>DA_FROM</type>
<position>52.5,-34</position>
<input>
<ID>IN_0</ID>545 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_bus</lparam></gate>
<gate>
<ID>45</ID>
<type>AI_REGISTER12</type>
<position>89,-46.5</position>
<input>
<ID>IN_0</ID>307 </input>
<input>
<ID>IN_1</ID>308 </input>
<input>
<ID>IN_10</ID>316 </input>
<input>
<ID>IN_11</ID>317 </input>
<input>
<ID>IN_2</ID>306 </input>
<input>
<ID>IN_3</ID>309 </input>
<input>
<ID>IN_4</ID>310 </input>
<input>
<ID>IN_5</ID>311 </input>
<input>
<ID>IN_6</ID>312 </input>
<input>
<ID>IN_7</ID>313 </input>
<input>
<ID>IN_8</ID>314 </input>
<input>
<ID>IN_9</ID>315 </input>
<output>
<ID>OUT_0</ID>384 </output>
<output>
<ID>OUT_1</ID>382 </output>
<output>
<ID>OUT_10</ID>385 </output>
<output>
<ID>OUT_11</ID>386 </output>
<output>
<ID>OUT_2</ID>388 </output>
<output>
<ID>OUT_3</ID>387 </output>
<output>
<ID>OUT_4</ID>378 </output>
<output>
<ID>OUT_5</ID>381 </output>
<output>
<ID>OUT_6</ID>379 </output>
<output>
<ID>OUT_7</ID>383 </output>
<output>
<ID>OUT_8</ID>389 </output>
<output>
<ID>OUT_9</ID>380 </output>
<input>
<ID>clear</ID>597 </input>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>count_enable</ID>596 </input>
<input>
<ID>load</ID>595 </input>
<gparam>VALUE_BOX -2.4,-0.8,2.4,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 12</lparam>
<lparam>MAX_COUNT 4095</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>239</ID>
<type>DA_FROM</type>
<position>96.5,-67.5</position>
<input>
<ID>IN_0</ID>591 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_LD</lparam></gate>
<gate>
<ID>47</ID>
<type>AM_REGISTER16</type>
<position>99.5,-78.5</position>
<input>
<ID>IN_0</ID>968 </input>
<input>
<ID>IN_1</ID>984 </input>
<input>
<ID>IN_10</ID>971 </input>
<input>
<ID>IN_11</ID>987 </input>
<input>
<ID>IN_12</ID>973 </input>
<input>
<ID>IN_13</ID>988 </input>
<input>
<ID>IN_14</ID>975 </input>
<input>
<ID>IN_15</ID>991 </input>
<input>
<ID>IN_2</ID>969 </input>
<input>
<ID>IN_3</ID>985 </input>
<input>
<ID>IN_4</ID>972 </input>
<input>
<ID>IN_5</ID>989 </input>
<input>
<ID>IN_6</ID>974 </input>
<input>
<ID>IN_7</ID>990 </input>
<input>
<ID>IN_8</ID>970 </input>
<input>
<ID>IN_9</ID>986 </input>
<output>
<ID>OUT_0</ID>563 </output>
<output>
<ID>OUT_1</ID>564 </output>
<output>
<ID>OUT_10</ID>573 </output>
<output>
<ID>OUT_11</ID>574 </output>
<output>
<ID>OUT_12</ID>575 </output>
<output>
<ID>OUT_13</ID>576 </output>
<output>
<ID>OUT_14</ID>577 </output>
<output>
<ID>OUT_15</ID>578 </output>
<output>
<ID>OUT_2</ID>565 </output>
<output>
<ID>OUT_3</ID>566 </output>
<output>
<ID>OUT_4</ID>567 </output>
<output>
<ID>OUT_5</ID>568 </output>
<output>
<ID>OUT_6</ID>569 </output>
<output>
<ID>OUT_7</ID>570 </output>
<output>
<ID>OUT_8</ID>571 </output>
<output>
<ID>OUT_9</ID>572 </output>
<input>
<ID>clear</ID>593 </input>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>count_enable</ID>592 </input>
<input>
<ID>load</ID>591 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>52</ID>
<type>BX_16X1_BUS_END</type>
<position>130.5,-44.5</position>
<input>
<ID>Bus_in_0</ID>362 </input>
<input>
<ID>IN_1</ID>363 </input>
<input>
<ID>IN_10</ID>377 </input>
<input>
<ID>IN_11</ID>371 </input>
<input>
<ID>IN_12</ID>372 </input>
<input>
<ID>IN_13</ID>375 </input>
<input>
<ID>IN_14</ID>376 </input>
<input>
<ID>IN_15</ID>374 </input>
<input>
<ID>IN_2</ID>368 </input>
<input>
<ID>IN_3</ID>364 </input>
<input>
<ID>IN_4</ID>365 </input>
<input>
<ID>IN_5</ID>366 </input>
<input>
<ID>IN_6</ID>369 </input>
<input>
<ID>IN_7</ID>367 </input>
<input>
<ID>IN_8</ID>370 </input>
<input>
<ID>IN_9</ID>373 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>116</ID>
<type>AE_REGISTER8</type>
<position>87.5,-147</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>198 </input>
<input>
<ID>IN_2</ID>199 </input>
<input>
<ID>IN_3</ID>196 </input>
<input>
<ID>IN_4</ID>197 </input>
<input>
<ID>IN_5</ID>200 </input>
<input>
<ID>IN_6</ID>194 </input>
<input>
<ID>IN_7</ID>201 </input>
<output>
<ID>OUT_0</ID>514 </output>
<output>
<ID>OUT_1</ID>518 </output>
<output>
<ID>OUT_2</ID>515 </output>
<output>
<ID>OUT_3</ID>516 </output>
<output>
<ID>OUT_4</ID>521 </output>
<output>
<ID>OUT_5</ID>519 </output>
<output>
<ID>OUT_6</ID>517 </output>
<output>
<ID>OUT_7</ID>520 </output>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>load</ID>202 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>270</ID>
<type>DA_FROM</type>
<position>87.5,-13.5</position>
<input>
<ID>IN_0</ID>708 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Mem_R</lparam></gate>
<gate>
<ID>245</ID>
<type>DA_FROM</type>
<position>116,-68</position>
<input>
<ID>IN_0</ID>594 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_bus</lparam></gate>
<gate>
<ID>53</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>119.5,-44.5</position>
<input>
<ID>ENABLE_0</ID>546 </input>
<input>
<ID>IN_0</ID>384 </input>
<input>
<ID>IN_1</ID>382 </input>
<input>
<ID>IN_10</ID>385 </input>
<input>
<ID>IN_11</ID>386 </input>
<input>
<ID>IN_2</ID>388 </input>
<input>
<ID>IN_3</ID>387 </input>
<input>
<ID>IN_4</ID>378 </input>
<input>
<ID>IN_5</ID>381 </input>
<input>
<ID>IN_6</ID>379 </input>
<input>
<ID>IN_7</ID>383 </input>
<input>
<ID>IN_8</ID>389 </input>
<input>
<ID>IN_9</ID>380 </input>
<output>
<ID>OUT_0</ID>362 </output>
<output>
<ID>OUT_1</ID>363 </output>
<output>
<ID>OUT_10</ID>377 </output>
<output>
<ID>OUT_11</ID>371 </output>
<output>
<ID>OUT_12</ID>372 </output>
<output>
<ID>OUT_13</ID>375 </output>
<output>
<ID>OUT_14</ID>376 </output>
<output>
<ID>OUT_15</ID>374 </output>
<output>
<ID>OUT_2</ID>368 </output>
<output>
<ID>OUT_3</ID>364 </output>
<output>
<ID>OUT_4</ID>365 </output>
<output>
<ID>OUT_5</ID>366 </output>
<output>
<ID>OUT_6</ID>369 </output>
<output>
<ID>OUT_7</ID>367 </output>
<output>
<ID>OUT_8</ID>370 </output>
<output>
<ID>OUT_9</ID>373 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>54</ID>
<type>BX_16X1_BUS_END</type>
<position>130.5,-78.5</position>
<input>
<ID>Bus_in_0</ID>390 </input>
<input>
<ID>IN_1</ID>391 </input>
<input>
<ID>IN_10</ID>405 </input>
<input>
<ID>IN_11</ID>399 </input>
<input>
<ID>IN_12</ID>400 </input>
<input>
<ID>IN_13</ID>403 </input>
<input>
<ID>IN_14</ID>404 </input>
<input>
<ID>IN_15</ID>402 </input>
<input>
<ID>IN_2</ID>396 </input>
<input>
<ID>IN_3</ID>392 </input>
<input>
<ID>IN_4</ID>393 </input>
<input>
<ID>IN_5</ID>394 </input>
<input>
<ID>IN_6</ID>397 </input>
<input>
<ID>IN_7</ID>395 </input>
<input>
<ID>IN_8</ID>398 </input>
<input>
<ID>IN_9</ID>401 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>247</ID>
<type>DA_FROM</type>
<position>86,-34.5</position>
<input>
<ID>IN_0</ID>595 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_LD</lparam></gate>
<gate>
<ID>1091</ID>
<type>DA_FROM</type>
<position>-60,-114</position>
<input>
<ID>IN_0</ID>1214 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>55</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>119.5,-78.5</position>
<input>
<ID>ENABLE_0</ID>594 </input>
<input>
<ID>IN_0</ID>563 </input>
<input>
<ID>IN_1</ID>564 </input>
<input>
<ID>IN_10</ID>573 </input>
<input>
<ID>IN_11</ID>574 </input>
<input>
<ID>IN_12</ID>575 </input>
<input>
<ID>IN_13</ID>576 </input>
<input>
<ID>IN_14</ID>577 </input>
<input>
<ID>IN_15</ID>578 </input>
<input>
<ID>IN_2</ID>565 </input>
<input>
<ID>IN_3</ID>566 </input>
<input>
<ID>IN_4</ID>567 </input>
<input>
<ID>IN_5</ID>568 </input>
<input>
<ID>IN_6</ID>569 </input>
<input>
<ID>IN_7</ID>570 </input>
<input>
<ID>IN_8</ID>571 </input>
<input>
<ID>IN_9</ID>572 </input>
<output>
<ID>OUT_0</ID>390 </output>
<output>
<ID>OUT_1</ID>391 </output>
<output>
<ID>OUT_10</ID>405 </output>
<output>
<ID>OUT_11</ID>399 </output>
<output>
<ID>OUT_12</ID>400 </output>
<output>
<ID>OUT_13</ID>403 </output>
<output>
<ID>OUT_14</ID>404 </output>
<output>
<ID>OUT_15</ID>402 </output>
<output>
<ID>OUT_2</ID>396 </output>
<output>
<ID>OUT_3</ID>392 </output>
<output>
<ID>OUT_4</ID>393 </output>
<output>
<ID>OUT_5</ID>394 </output>
<output>
<ID>OUT_6</ID>397 </output>
<output>
<ID>OUT_7</ID>395 </output>
<output>
<ID>OUT_8</ID>398 </output>
<output>
<ID>OUT_9</ID>401 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>231</ID>
<type>DA_FROM</type>
<position>86,-132</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_CLR</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>-49,-57.5</position>
<output>
<ID>OUT_0</ID>488 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>312</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>148.5,-57.5</position>
<input>
<ID>IN_0</ID>843 </input>
<input>
<ID>IN_1</ID>864 </input>
<input>
<ID>IN_2</ID>844 </input>
<input>
<ID>IN_3</ID>863 </input>
<input>
<ID>IN_4</ID>865 </input>
<input>
<ID>IN_5</ID>839 </input>
<input>
<ID>IN_6</ID>869 </input>
<input>
<ID>IN_7</ID>870 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>167</ID>
<type>DA_FROM</type>
<position>22.5,-57</position>
<input>
<ID>IN_0</ID>544 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_CLR</lparam></gate>
<gate>
<ID>251</ID>
<type>DA_FROM</type>
<position>86,-57</position>
<input>
<ID>IN_0</ID>597 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_CLR</lparam></gate>
<gate>
<ID>123</ID>
<type>DA_FROM</type>
<position>3.5,-55</position>
<input>
<ID>IN_0</ID>513 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_LABEL</type>
<position>-3.5,-44</position>
<gparam>LABEL_TEXT Address Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>146,-78</position>
<gparam>LABEL_TEXT Accumulator</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>AA_LABEL</type>
<position>-1,-78</position>
<gparam>LABEL_TEXT Data Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>131</ID>
<type>AA_LABEL</type>
<position>-6.5,-119</position>
<gparam>LABEL_TEXT Instruction Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>AA_LABEL</type>
<position>149.5,-44</position>
<gparam>LABEL_TEXT Program Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_LABEL</type>
<position>147.5,-118.5</position>
<gparam>LABEL_TEXT Temp Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>137</ID>
<type>AA_LABEL</type>
<position>116,-146</position>
<gparam>LABEL_TEXT Output Register</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>98,-147</position>
<input>
<ID>IN_0</ID>514 </input>
<input>
<ID>IN_1</ID>518 </input>
<input>
<ID>IN_2</ID>515 </input>
<input>
<ID>IN_3</ID>516 </input>
<input>
<ID>IN_4</ID>521 </input>
<input>
<ID>IN_5</ID>519 </input>
<input>
<ID>IN_6</ID>517 </input>
<input>
<ID>IN_7</ID>520 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>1055</ID>
<type>AA_LABEL</type>
<position>-49,-34.5</position>
<gparam>LABEL_TEXT Turn switch on for one or two</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>116,-34</position>
<input>
<ID>IN_0</ID>546 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_bus</lparam></gate>
<gate>
<ID>217</ID>
<type>DA_FROM</type>
<position>22.5,-67.5</position>
<input>
<ID>IN_0</ID>580 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_LD</lparam></gate>
<gate>
<ID>219</ID>
<type>DA_FROM</type>
<position>22.5,-65</position>
<input>
<ID>IN_0</ID>581 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_INC</lparam></gate>
<gate>
<ID>241</ID>
<type>DA_FROM</type>
<position>96.5,-64.5</position>
<input>
<ID>IN_0</ID>592 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_INC</lparam></gate>
<gate>
<ID>243</ID>
<type>DA_FROM</type>
<position>96.5,-91</position>
<input>
<ID>IN_0</ID>593 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_CLR</lparam></gate>
<gate>
<ID>249</ID>
<type>DA_FROM</type>
<position>86,-32</position>
<input>
<ID>IN_0</ID>596 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_INC</lparam></gate>
<gate>
<ID>6</ID>
<type>BX_16X1_BUS_END</type>
<position>74,-26</position>
<input>
<ID>Bus_in_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<input>
<ID>IN_10</ID>68 </input>
<input>
<ID>IN_11</ID>69 </input>
<input>
<ID>IN_12</ID>60 </input>
<input>
<ID>IN_13</ID>62 </input>
<input>
<ID>IN_14</ID>72 </input>
<input>
<ID>IN_15</ID>70 </input>
<input>
<ID>IN_2</ID>57 </input>
<input>
<ID>IN_3</ID>63 </input>
<input>
<ID>IN_4</ID>64 </input>
<input>
<ID>IN_5</ID>61 </input>
<input>
<ID>IN_6</ID>65 </input>
<input>
<ID>IN_7</ID>66 </input>
<input>
<ID>IN_8</ID>71 </input>
<input>
<ID>IN_9</ID>67 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>860</ID>
<type>DA_FROM</type>
<position>82.5,-77</position>
<input>
<ID>IN_0</ID>986 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi9</lparam></gate>
<gate>
<ID>13</ID>
<type>AM_REGISTER16</type>
<position>89,-119.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>139 </input>
<input>
<ID>IN_10</ID>153 </input>
<input>
<ID>IN_11</ID>141 </input>
<input>
<ID>IN_12</ID>142 </input>
<input>
<ID>IN_13</ID>154 </input>
<input>
<ID>IN_14</ID>147 </input>
<input>
<ID>IN_15</ID>143 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>140 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>151 </input>
<input>
<ID>IN_6</ID>145 </input>
<input>
<ID>IN_7</ID>152 </input>
<input>
<ID>IN_8</ID>144 </input>
<input>
<ID>IN_9</ID>146 </input>
<output>
<ID>OUT_0</ID>182 </output>
<output>
<ID>OUT_1</ID>155 </output>
<output>
<ID>OUT_10</ID>180 </output>
<output>
<ID>OUT_11</ID>181 </output>
<output>
<ID>OUT_12</ID>183 </output>
<output>
<ID>OUT_13</ID>185 </output>
<output>
<ID>OUT_14</ID>184 </output>
<output>
<ID>OUT_15</ID>74 </output>
<output>
<ID>OUT_2</ID>156 </output>
<output>
<ID>OUT_3</ID>157 </output>
<output>
<ID>OUT_4</ID>158 </output>
<output>
<ID>OUT_5</ID>159 </output>
<output>
<ID>OUT_6</ID>160 </output>
<output>
<ID>OUT_7</ID>161 </output>
<output>
<ID>OUT_8</ID>178 </output>
<output>
<ID>OUT_9</ID>179 </output>
<input>
<ID>clear</ID>190 </input>
<input>
<ID>clock</ID>513 </input>
<input>
<ID>count_enable</ID>188 </input>
<input>
<ID>load</ID>187 </input>
<gparam>VALUE_BOX -2.8,-0.8,2.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 16</lparam>
<lparam>MAX_COUNT 65536</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>14</ID>
<type>BX_16X1_BUS_END</type>
<position>130.5,-119.5</position>
<input>
<ID>Bus_in_0</ID>91 </input>
<input>
<ID>IN_1</ID>92 </input>
<input>
<ID>IN_10</ID>138 </input>
<input>
<ID>IN_11</ID>132 </input>
<input>
<ID>IN_12</ID>133 </input>
<input>
<ID>IN_13</ID>136 </input>
<input>
<ID>IN_14</ID>137 </input>
<input>
<ID>IN_15</ID>73 </input>
<input>
<ID>IN_2</ID>113 </input>
<input>
<ID>IN_3</ID>93 </input>
<input>
<ID>IN_4</ID>94 </input>
<input>
<ID>IN_5</ID>95 </input>
<input>
<ID>IN_6</ID>130 </input>
<input>
<ID>IN_7</ID>96 </input>
<input>
<ID>IN_8</ID>131 </input>
<input>
<ID>IN_9</ID>134 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>15</ID>
<type>BU_TRI_STATE_16BIT</type>
<position>119.5,-119.5</position>
<input>
<ID>ENABLE_0</ID>193 </input>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>155 </input>
<input>
<ID>IN_10</ID>180 </input>
<input>
<ID>IN_11</ID>181 </input>
<input>
<ID>IN_12</ID>183 </input>
<input>
<ID>IN_13</ID>185 </input>
<input>
<ID>IN_14</ID>184 </input>
<input>
<ID>IN_15</ID>74 </input>
<input>
<ID>IN_2</ID>156 </input>
<input>
<ID>IN_3</ID>157 </input>
<input>
<ID>IN_4</ID>158 </input>
<input>
<ID>IN_5</ID>159 </input>
<input>
<ID>IN_6</ID>160 </input>
<input>
<ID>IN_7</ID>161 </input>
<input>
<ID>IN_8</ID>178 </input>
<input>
<ID>IN_9</ID>179 </input>
<output>
<ID>OUT_0</ID>91 </output>
<output>
<ID>OUT_1</ID>92 </output>
<output>
<ID>OUT_10</ID>138 </output>
<output>
<ID>OUT_11</ID>132 </output>
<output>
<ID>OUT_12</ID>133 </output>
<output>
<ID>OUT_13</ID>136 </output>
<output>
<ID>OUT_14</ID>137 </output>
<output>
<ID>OUT_15</ID>73 </output>
<output>
<ID>OUT_2</ID>113 </output>
<output>
<ID>OUT_3</ID>93 </output>
<output>
<ID>OUT_4</ID>94 </output>
<output>
<ID>OUT_5</ID>95 </output>
<output>
<ID>OUT_6</ID>130 </output>
<output>
<ID>OUT_7</ID>96 </output>
<output>
<ID>OUT_8</ID>131 </output>
<output>
<ID>OUT_9</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>864</ID>
<type>DA_FROM</type>
<position>82.5,-73</position>
<input>
<ID>IN_0</ID>988 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi13</lparam></gate>
<gate>
<ID>17</ID>
<type>BX_16X1_BUS_END</type>
<position>81,-119.5</position>
<input>
<ID>Bus_in_0</ID>150 </input>
<input>
<ID>IN_1</ID>139 </input>
<input>
<ID>IN_10</ID>153 </input>
<input>
<ID>IN_11</ID>141 </input>
<input>
<ID>IN_12</ID>142 </input>
<input>
<ID>IN_13</ID>154 </input>
<input>
<ID>IN_14</ID>147 </input>
<input>
<ID>IN_15</ID>143 </input>
<input>
<ID>IN_2</ID>149 </input>
<input>
<ID>IN_3</ID>140 </input>
<input>
<ID>IN_4</ID>148 </input>
<input>
<ID>IN_5</ID>151 </input>
<input>
<ID>IN_6</ID>145 </input>
<input>
<ID>IN_7</ID>152 </input>
<input>
<ID>IN_8</ID>144 </input>
<input>
<ID>IN_9</ID>146 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>24</ID>
<type>DA_FROM</type>
<position>52.5,-109</position>
<input>
<ID>IN_0</ID>192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR_bus</lparam></gate>
<gate>
<ID>26</ID>
<type>DA_FROM</type>
<position>116,-109</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_bus</lparam></gate>
<gate>
<ID>28</ID>
<type>BX_16X1_BUS_END</type>
<position>80.5,-142.5</position>
<input>
<ID>Bus_in_0</ID>195 </input>
<input>
<ID>IN_1</ID>198 </input>
<input>
<ID>IN_2</ID>199 </input>
<input>
<ID>IN_3</ID>196 </input>
<input>
<ID>IN_4</ID>197 </input>
<input>
<ID>IN_5</ID>200 </input>
<input>
<ID>IN_6</ID>194 </input>
<input>
<ID>IN_7</ID>201 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>34</ID>
<type>DA_FROM</type>
<position>89.5,-138.5</position>
<input>
<ID>IN_0</ID>202 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID OUTR_LD</lparam></gate>
<gate>
<ID>4</ID>
<type>DE_TO</type>
<position>116,-90.5</position>
<input>
<ID>IN_0</ID>563 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>11</ID>
<type>DE_TO</type>
<position>125.5,-91.5</position>
<input>
<ID>IN_0</ID>564 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo1</lparam></gate>
<gate>
<ID>12</ID>
<type>DE_TO</type>
<position>116,-92.5</position>
<input>
<ID>IN_0</ID>565 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo2</lparam></gate>
<gate>
<ID>19</ID>
<type>DE_TO</type>
<position>125.5,-93.5</position>
<input>
<ID>IN_0</ID>566 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo3</lparam></gate>
<gate>
<ID>21</ID>
<type>DE_TO</type>
<position>116,-94.5</position>
<input>
<ID>IN_0</ID>567 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo4</lparam></gate>
<gate>
<ID>23</ID>
<type>DE_TO</type>
<position>125.5,-95.5</position>
<input>
<ID>IN_0</ID>568 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo5</lparam></gate>
<gate>
<ID>25</ID>
<type>DE_TO</type>
<position>116,-96.5</position>
<input>
<ID>IN_0</ID>569 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo6</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>125.5,-97.5</position>
<input>
<ID>IN_0</ID>570 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo7</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>116,-98.5</position>
<input>
<ID>IN_0</ID>571 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo8</lparam></gate>
<gate>
<ID>33</ID>
<type>DE_TO</type>
<position>125.5,-99.5</position>
<input>
<ID>IN_0</ID>572 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo9</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>116,-100.5</position>
<input>
<ID>IN_0</ID>573 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo10</lparam></gate>
<gate>
<ID>38</ID>
<type>DE_TO</type>
<position>125.5,-101.5</position>
<input>
<ID>IN_0</ID>574 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo11</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>116,-102.5</position>
<input>
<ID>IN_0</ID>575 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo12</lparam></gate>
<gate>
<ID>1094</ID>
<type>DE_TO</type>
<position>-50,-106</position>
<input>
<ID>IN_0</ID>1215 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR0</lparam></gate>
<gate>
<ID>42</ID>
<type>DE_TO</type>
<position>125.5,-103.5</position>
<input>
<ID>IN_0</ID>576 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo13</lparam></gate>
<gate>
<ID>43</ID>
<type>DE_TO</type>
<position>116,-104.5</position>
<input>
<ID>IN_0</ID>577 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo14</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>125.5,-105.5</position>
<input>
<ID>IN_0</ID>578 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>71</ID>
<type>DE_TO</type>
<position>20.5,-17.5</position>
<input>
<ID>IN_0</ID>1 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR0</lparam></gate>
<gate>
<ID>72</ID>
<type>DE_TO</type>
<position>28.5,-16.5</position>
<input>
<ID>IN_0</ID>12 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR1</lparam></gate>
<gate>
<ID>73</ID>
<type>DE_TO</type>
<position>20.5,-15.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR2</lparam></gate>
<gate>
<ID>74</ID>
<type>DE_TO</type>
<position>28.5,-14.5</position>
<input>
<ID>IN_0</ID>10 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR3</lparam></gate>
<gate>
<ID>1087</ID>
<type>AE_REGISTER8</type>
<position>-57,-103</position>
<input>
<ID>IN_0</ID>1213 </input>
<input>
<ID>IN_1</ID>1212 </input>
<input>
<ID>IN_2</ID>1211 </input>
<input>
<ID>IN_3</ID>1210 </input>
<input>
<ID>IN_4</ID>1206 </input>
<input>
<ID>IN_5</ID>1207 </input>
<input>
<ID>IN_6</ID>1208 </input>
<input>
<ID>IN_7</ID>1209 </input>
<output>
<ID>OUT_0</ID>1215 </output>
<output>
<ID>OUT_1</ID>1219 </output>
<output>
<ID>OUT_2</ID>1218 </output>
<output>
<ID>OUT_3</ID>1220 </output>
<output>
<ID>OUT_4</ID>1216 </output>
<output>
<ID>OUT_5</ID>1222 </output>
<output>
<ID>OUT_6</ID>1217 </output>
<output>
<ID>OUT_7</ID>1221 </output>
<input>
<ID>clock</ID>1214 </input>
<input>
<ID>load</ID>1223 </input>
<gparam>VALUE_BOX -1.8,-0.8,1.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>MAX_COUNT 255</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>75</ID>
<type>DE_TO</type>
<position>20.5,-13.5</position>
<input>
<ID>IN_0</ID>9 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR4</lparam></gate>
<gate>
<ID>76</ID>
<type>DE_TO</type>
<position>28.5,-12.5</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR5</lparam></gate>
<gate>
<ID>77</ID>
<type>DE_TO</type>
<position>20.5,-11.5</position>
<input>
<ID>IN_0</ID>7 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR6</lparam></gate>
<gate>
<ID>1074</ID>
<type>AA_LABEL</type>
<position>-48.5,-38.5</position>
<gparam>LABEL_TEXT Then switch back off to start the</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>DE_TO</type>
<position>28.5,-10.5</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR7</lparam></gate>
<gate>
<ID>79</ID>
<type>DE_TO</type>
<position>20.5,-9.5</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR8</lparam></gate>
<gate>
<ID>80</ID>
<type>DE_TO</type>
<position>28.5,-8.5</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR9</lparam></gate>
<gate>
<ID>81</ID>
<type>DE_TO</type>
<position>20.5,-7.5</position>
<input>
<ID>IN_0</ID>3 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR10</lparam></gate>
<gate>
<ID>82</ID>
<type>DE_TO</type>
<position>28.5,-6.5</position>
<input>
<ID>IN_0</ID>2 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID AR11</lparam></gate>
<gate>
<ID>84</ID>
<type>DE_TO</type>
<position>42,-91</position>
<input>
<ID>IN_0</ID>547 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR0</lparam></gate>
<gate>
<ID>1081</ID>
<type>DE_TO</type>
<position>-52.5,-74.5</position>
<input>
<ID>IN_0</ID>1204 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI_SET</lparam></gate>
<gate>
<ID>85</ID>
<type>DE_TO</type>
<position>50.5,-92</position>
<input>
<ID>IN_0</ID>548 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR1</lparam></gate>
<gate>
<ID>1082</ID>
<type>DE_TO</type>
<position>-52.5,-78.5</position>
<input>
<ID>IN_0</ID>1205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO_SET</lparam></gate>
<gate>
<ID>86</ID>
<type>DE_TO</type>
<position>42,-93</position>
<input>
<ID>IN_0</ID>549 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR2</lparam></gate>
<gate>
<ID>87</ID>
<type>DE_TO</type>
<position>50.5,-94</position>
<input>
<ID>IN_0</ID>550 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR3</lparam></gate>
<gate>
<ID>88</ID>
<type>DE_TO</type>
<position>42,-95</position>
<input>
<ID>IN_0</ID>551 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR4</lparam></gate>
<gate>
<ID>89</ID>
<type>DE_TO</type>
<position>50.5,-96</position>
<input>
<ID>IN_0</ID>552 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR5</lparam></gate>
<gate>
<ID>91</ID>
<type>DE_TO</type>
<position>42,-97</position>
<input>
<ID>IN_0</ID>553 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR6</lparam></gate>
<gate>
<ID>92</ID>
<type>DE_TO</type>
<position>50.5,-98</position>
<input>
<ID>IN_0</ID>554 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR7</lparam></gate>
<gate>
<ID>93</ID>
<type>DE_TO</type>
<position>42,-99</position>
<input>
<ID>IN_0</ID>555 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR8</lparam></gate>
<gate>
<ID>94</ID>
<type>DE_TO</type>
<position>50.5,-100</position>
<input>
<ID>IN_0</ID>556 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR9</lparam></gate>
<gate>
<ID>95</ID>
<type>DE_TO</type>
<position>42,-101</position>
<input>
<ID>IN_0</ID>557 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR10</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>50.5,-102</position>
<input>
<ID>IN_0</ID>558 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR11</lparam></gate>
<gate>
<ID>98</ID>
<type>DE_TO</type>
<position>42,-103</position>
<input>
<ID>IN_0</ID>559 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR12</lparam></gate>
<gate>
<ID>100</ID>
<type>DE_TO</type>
<position>50.5,-104</position>
<input>
<ID>IN_0</ID>560 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR13</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>42,-105</position>
<input>
<ID>IN_0</ID>561 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR14</lparam></gate>
<gate>
<ID>104</ID>
<type>DE_TO</type>
<position>50.5,-106</position>
<input>
<ID>IN_0</ID>562 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR15</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>42,-132</position>
<input>
<ID>IN_0</ID>285 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR0</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>50.5,-133</position>
<input>
<ID>IN_0</ID>274 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR1</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>42,-134</position>
<input>
<ID>IN_0</ID>275 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR2</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>50.5,-135</position>
<input>
<ID>IN_0</ID>276 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR3</lparam></gate>
<gate>
<ID>111</ID>
<type>DE_TO</type>
<position>42,-136</position>
<input>
<ID>IN_0</ID>277 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR4</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>50.5,-137</position>
<input>
<ID>IN_0</ID>278 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR5</lparam></gate>
<gate>
<ID>113</ID>
<type>DE_TO</type>
<position>42,-138</position>
<input>
<ID>IN_0</ID>279 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR6</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>50.5,-139</position>
<input>
<ID>IN_0</ID>280 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR7</lparam></gate>
<gate>
<ID>115</ID>
<type>DE_TO</type>
<position>42,-140</position>
<input>
<ID>IN_0</ID>281 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR8</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>50.5,-141</position>
<input>
<ID>IN_0</ID>282 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR9</lparam></gate>
<gate>
<ID>118</ID>
<type>DE_TO</type>
<position>42,-142</position>
<input>
<ID>IN_0</ID>283 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR10</lparam></gate>
<gate>
<ID>119</ID>
<type>DE_TO</type>
<position>50.5,-143</position>
<input>
<ID>IN_0</ID>284 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR11</lparam></gate>
<gate>
<ID>120</ID>
<type>DE_TO</type>
<position>42,-144</position>
<input>
<ID>IN_0</ID>286 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR12</lparam></gate>
<gate>
<ID>121</ID>
<type>DE_TO</type>
<position>50.5,-145</position>
<input>
<ID>IN_0</ID>288 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR13</lparam></gate>
<gate>
<ID>122</ID>
<type>DE_TO</type>
<position>42,-146</position>
<input>
<ID>IN_0</ID>287 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR14</lparam></gate>
<gate>
<ID>124</ID>
<type>DE_TO</type>
<position>50.5,-147</position>
<input>
<ID>IN_0</ID>289 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR15</lparam></gate>
<gate>
<ID>267</ID>
<type>DA_FROM</type>
<position>87.5,-11.5</position>
<input>
<ID>IN_0</ID>662 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Mem_W</lparam></gate>
<gate>
<ID>304</ID>
<type>BX_16X1_BUS_END</type>
<position>139.5,-61.5</position>
<input>
<ID>Bus_in_0</ID>811 </input>
<input>
<ID>IN_1</ID>837 </input>
<input>
<ID>IN_10</ID>844 </input>
<input>
<ID>IN_11</ID>863 </input>
<input>
<ID>IN_12</ID>865 </input>
<input>
<ID>IN_13</ID>839 </input>
<input>
<ID>IN_14</ID>869 </input>
<input>
<ID>IN_15</ID>870 </input>
<input>
<ID>IN_2</ID>817 </input>
<input>
<ID>IN_3</ID>838 </input>
<input>
<ID>IN_4</ID>813 </input>
<input>
<ID>IN_5</ID>792 </input>
<input>
<ID>IN_6</ID>818 </input>
<input>
<ID>IN_7</ID>812 </input>
<input>
<ID>IN_8</ID>843 </input>
<input>
<ID>IN_9</ID>864 </input>
<input>
<ID>OUT</ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </input>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 16</lparam></gate>
<gate>
<ID>310</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>148.5,-66.5</position>
<input>
<ID>IN_0</ID>811 </input>
<input>
<ID>IN_1</ID>837 </input>
<input>
<ID>IN_2</ID>817 </input>
<input>
<ID>IN_3</ID>838 </input>
<input>
<ID>IN_4</ID>813 </input>
<input>
<ID>IN_5</ID>792 </input>
<input>
<ID>IN_6</ID>818 </input>
<input>
<ID>IN_7</ID>812 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>851</ID>
<type>DA_FROM</type>
<position>91.5,-86</position>
<input>
<ID>IN_0</ID>968 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi0</lparam></gate>
<gate>
<ID>852</ID>
<type>DA_FROM</type>
<position>82.5,-85</position>
<input>
<ID>IN_0</ID>984 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi1</lparam></gate>
<gate>
<ID>853</ID>
<type>DA_FROM</type>
<position>91.5,-84</position>
<input>
<ID>IN_0</ID>969 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi2</lparam></gate>
<gate>
<ID>854</ID>
<type>DA_FROM</type>
<position>82.5,-83</position>
<input>
<ID>IN_0</ID>985 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi3</lparam></gate>
<gate>
<ID>855</ID>
<type>DA_FROM</type>
<position>91.5,-82</position>
<input>
<ID>IN_0</ID>972 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi4</lparam></gate>
<gate>
<ID>856</ID>
<type>DA_FROM</type>
<position>82.5,-81</position>
<input>
<ID>IN_0</ID>989 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi5</lparam></gate>
<gate>
<ID>857</ID>
<type>DA_FROM</type>
<position>91.5,-80</position>
<input>
<ID>IN_0</ID>974 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi6</lparam></gate>
<gate>
<ID>858</ID>
<type>DA_FROM</type>
<position>82.5,-79</position>
<input>
<ID>IN_0</ID>990 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi7</lparam></gate>
<gate>
<ID>859</ID>
<type>DA_FROM</type>
<position>91.5,-78</position>
<input>
<ID>IN_0</ID>970 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi8</lparam></gate>
<gate>
<ID>861</ID>
<type>DA_FROM</type>
<position>91.5,-76</position>
<input>
<ID>IN_0</ID>971 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi10</lparam></gate>
<gate>
<ID>862</ID>
<type>DA_FROM</type>
<position>82.5,-75</position>
<input>
<ID>IN_0</ID>987 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi11</lparam></gate>
<gate>
<ID>863</ID>
<type>DA_FROM</type>
<position>91.5,-74</position>
<input>
<ID>IN_0</ID>973 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi12</lparam></gate>
<gate>
<ID>865</ID>
<type>DA_FROM</type>
<position>91.5,-72</position>
<input>
<ID>IN_0</ID>975 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi14</lparam></gate>
<gate>
<ID>866</ID>
<type>DA_FROM</type>
<position>82.5,-71</position>
<input>
<ID>IN_0</ID>991 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi15</lparam></gate>
<gate>
<ID>1089</ID>
<type>DE_TO</type>
<position>-50,-104</position>
<input>
<ID>IN_0</ID>1218 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR2</lparam></gate>
<gate>
<ID>221</ID>
<type>DA_FROM</type>
<position>22.5,-91</position>
<input>
<ID>IN_0</ID>582 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_CLR</lparam></gate>
<gate>
<ID>547</ID>
<type>AA_TOGGLE</type>
<position>-54.5,-44.5</position>
<output>
<ID>OUT_0</ID>907 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>670</ID>
<type>DE_TO</type>
<position>-49,-44.5</position>
<input>
<ID>IN_0</ID>907 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>1036</ID>
<type>AA_LABEL</type>
<position>-49.5,-54.5</position>
<gparam>LABEL_TEXT Switch between manual and automatic clocking</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1046</ID>
<type>AA_LABEL</type>
<position>-49,-31.5</position>
<gparam>LABEL_TEXT START BUTTON</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1064</ID>
<type>AA_LABEL</type>
<position>-48,-36.5</position>
<gparam>LABEL_TEXT clock cycles to reset all the registers.</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1077</ID>
<type>AA_LABEL</type>
<position>-49,-40.5</position>
<gparam>LABEL_TEXT program loaded into memory</gparam>
<gparam>TEXT_HEIGHT 1.5</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1079</ID>
<type>AA_TOGGLE</type>
<position>-57.5,-74.5</position>
<output>
<ID>OUT_0</ID>1204 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1083</ID>
<type>AA_TOGGLE</type>
<position>-57.5,-78.5</position>
<output>
<ID>OUT_0</ID>1205 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1085</ID>
<type>AA_LABEL</type>
<position>-51,-71</position>
<gparam>LABEL_TEXT Set input and output flags</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1086</ID>
<type>DD_KEYPAD_HEX</type>
<position>-68.5,-96</position>
<output>
<ID>OUT_0</ID>1206 </output>
<output>
<ID>OUT_1</ID>1207 </output>
<output>
<ID>OUT_2</ID>1208 </output>
<output>
<ID>OUT_3</ID>1209 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1088</ID>
<type>DD_KEYPAD_HEX</type>
<position>-68.5,-109</position>
<output>
<ID>OUT_0</ID>1213 </output>
<output>
<ID>OUT_1</ID>1212 </output>
<output>
<ID>OUT_2</ID>1211 </output>
<output>
<ID>OUT_3</ID>1210 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1090</ID>
<type>DE_TO</type>
<position>-50,-100</position>
<input>
<ID>IN_0</ID>1217 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR6</lparam></gate>
<gate>
<ID>1095</ID>
<type>DE_TO</type>
<position>-41,-103</position>
<input>
<ID>IN_0</ID>1220 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR3</lparam></gate>
<gate>
<ID>1096</ID>
<type>DE_TO</type>
<position>-41,-101</position>
<input>
<ID>IN_0</ID>1222 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR5</lparam></gate>
<gate>
<ID>1098</ID>
<type>EE_VDD</type>
<position>-58,-95</position>
<output>
<ID>OUT_0</ID>1223 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>1099</ID>
<type>AA_LABEL</type>
<position>-51.5,-88</position>
<gparam>LABEL_TEXT Input register</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>41 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-52,65,-52</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<connection>
<GID>18</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>50 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-41,65,-41</points>
<connection>
<GID>20</GID>
<name>OUT_11</name></connection>
<connection>
<GID>18</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>544 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-57,26.5,-54</points>
<connection>
<GID>10</GID>
<name>clear</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-57,26.5,-57</points>
<connection>
<GID>167</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>401 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-77,128.5,-77</points>
<connection>
<GID>55</GID>
<name>OUT_9</name></connection>
<connection>
<GID>54</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-51,65,-51</points>
<connection>
<GID>20</GID>
<name>OUT_1</name></connection>
<connection>
<GID>18</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>56 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-42,65,-42</points>
<connection>
<GID>20</GID>
<name>OUT_10</name></connection>
<connection>
<GID>18</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-40,65,-40</points>
<connection>
<GID>20</GID>
<name>OUT_12</name></connection>
<connection>
<GID>18</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-39,65,-39</points>
<connection>
<GID>20</GID>
<name>OUT_13</name></connection>
<connection>
<GID>18</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>970 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-78,94.5,-78</points>
<connection>
<GID>47</GID>
<name>IN_8</name></connection>
<connection>
<GID>859</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1211 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-108,-62.5,-104</points>
<intersection>-108 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-108,-62.5,-108</points>
<connection>
<GID>1088</GID>
<name>OUT_2</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62.5,-104,-61,-104</points>
<connection>
<GID>1087</GID>
<name>IN_2</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-50,65,-50</points>
<connection>
<GID>20</GID>
<name>OUT_2</name></connection>
<connection>
<GID>18</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-38,65,-38</points>
<connection>
<GID>20</GID>
<name>OUT_14</name></connection>
<connection>
<GID>18</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-37,65,-37</points>
<connection>
<GID>20</GID>
<name>OUT_15</name></connection>
<connection>
<GID>18</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-49,65,-49</points>
<connection>
<GID>20</GID>
<name>OUT_3</name></connection>
<connection>
<GID>18</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-79,128.5,-79</points>
<connection>
<GID>55</GID>
<name>OUT_7</name></connection>
<connection>
<GID>54</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-48,65,-48</points>
<connection>
<GID>20</GID>
<name>OUT_4</name></connection>
<connection>
<GID>18</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-47,65,-47</points>
<connection>
<GID>20</GID>
<name>OUT_5</name></connection>
<connection>
<GID>18</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-46,65,-46</points>
<connection>
<GID>20</GID>
<name>OUT_6</name></connection>
<connection>
<GID>18</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>405 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-76,128.5,-76</points>
<connection>
<GID>55</GID>
<name>OUT_10</name></connection>
<connection>
<GID>54</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-45,65,-45</points>
<connection>
<GID>20</GID>
<name>OUT_7</name></connection>
<connection>
<GID>18</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>49 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-44,65,-44</points>
<connection>
<GID>20</GID>
<name>OUT_8</name></connection>
<connection>
<GID>18</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>403 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-73,128.5,-73</points>
<connection>
<GID>55</GID>
<name>OUT_13</name></connection>
<connection>
<GID>54</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-43,65,-43</points>
<connection>
<GID>20</GID>
<name>OUT_9</name></connection>
<connection>
<GID>18</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>378 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-48,117.5,-48</points>
<connection>
<GID>45</GID>
<name>OUT_4</name></connection>
<connection>
<GID>53</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>225 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-75,20.5,-75</points>
<connection>
<GID>40</GID>
<name>IN_11</name></connection>
<connection>
<GID>2</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>543 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-39,25.5,-32</points>
<connection>
<GID>10</GID>
<name>count_enable</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-32,25.5,-32</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1213 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-112,-61.5,-106</points>
<intersection>-112 1</intersection>
<intersection>-106 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-112,-61.5,-112</points>
<connection>
<GID>1088</GID>
<name>OUT_0</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-61.5,-106,-61,-106</points>
<connection>
<GID>1087</GID>
<name>IN_0</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-48,20.5,-48</points>
<connection>
<GID>16</GID>
<name>IN_4</name></connection>
<connection>
<GID>10</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>97 98 99 100 101 102 103 104 105 106 107 108 109 110 111 112 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-30,135,-30</points>
<intersection>13 10</intersection>
<intersection>74 44</intersection>
<intersection>135 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>135,-119.5,135,-30</points>
<intersection>-119.5 71</intersection>
<intersection>-78.5 35</intersection>
<intersection>-61.5 83</intersection>
<intersection>-44.5 32</intersection>
<intersection>-30 1</intersection></vsegment>
<vsegment>
<ID>10</ID>
<points>13,-119.5,13,-30</points>
<intersection>-119.5 81</intersection>
<intersection>-78.5 24</intersection>
<intersection>-44.5 14</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>13,-44.5,15.5,-44.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>13 10</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>13,-78.5,15.5,-78.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>13 10</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>132.5,-44.5,135,-44.5</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>135 4</intersection></hsegment>
<hsegment>
<ID>35</ID>
<points>132.5,-78.5,135,-78.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>135 4</intersection></hsegment>
<vsegment>
<ID>44</ID>
<points>74,-142.5,74,-28</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-142.5 77</intersection>
<intersection>-119.5 82</intersection>
<intersection>-78.5 50</intersection>
<intersection>-44.5 46</intersection>
<intersection>-30 1</intersection></vsegment>
<hsegment>
<ID>46</ID>
<points>69,-44.5,79,-44.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<intersection>74 44</intersection></hsegment>
<hsegment>
<ID>50</ID>
<points>69,-78.5,74,-78.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>74 44</intersection></hsegment>
<hsegment>
<ID>71</ID>
<points>132.5,-119.5,135,-119.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>135 4</intersection></hsegment>
<hsegment>
<ID>77</ID>
<points>74,-142.5,78.5,-142.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>74 44</intersection></hsegment>
<hsegment>
<ID>81</ID>
<points>13,-119.5,15.5,-119.5</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<intersection>13 10</intersection></hsegment>
<hsegment>
<ID>82</ID>
<points>69,-119.5,79,-119.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>74 44</intersection></hsegment>
<hsegment>
<ID>83</ID>
<points>135,-61.5,137.5,-61.5</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<intersection>135 4</intersection></hsegment></shape></wire>
<wire>
<ID>1214 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-114,-58,-108</points>
<connection>
<GID>1091</GID>
<name>IN_0</name></connection>
<connection>
<GID>1087</GID>
<name>clock</name></connection></vsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-82,128.5,-82</points>
<connection>
<GID>55</GID>
<name>OUT_4</name></connection>
<connection>
<GID>54</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-47,20.5,-47</points>
<connection>
<GID>16</GID>
<name>IN_5</name></connection>
<connection>
<GID>10</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-46,20.5,-46</points>
<connection>
<GID>16</GID>
<name>IN_6</name></connection>
<connection>
<GID>10</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>974 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-80,94.5,-80</points>
<connection>
<GID>47</GID>
<name>IN_6</name></connection>
<connection>
<GID>857</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-49,117.5,-49</points>
<connection>
<GID>45</GID>
<name>OUT_3</name></connection>
<connection>
<GID>53</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-45,20.5,-45</points>
<connection>
<GID>16</GID>
<name>IN_7</name></connection>
<connection>
<GID>10</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-44,20.5,-44</points>
<connection>
<GID>16</GID>
<name>IN_8</name></connection>
<connection>
<GID>10</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-80,128.5,-80</points>
<connection>
<GID>55</GID>
<name>OUT_6</name></connection>
<connection>
<GID>54</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-43,20.5,-43</points>
<connection>
<GID>16</GID>
<name>IN_9</name></connection>
<connection>
<GID>10</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-42,20.5,-42</points>
<connection>
<GID>16</GID>
<name>IN_10</name></connection>
<connection>
<GID>10</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-41,20.5,-41</points>
<connection>
<GID>16</GID>
<name>IN_11</name></connection>
<connection>
<GID>10</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-52,20.5,-52</points>
<connection>
<GID>16</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>10</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>374 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-37,128.5,-37</points>
<connection>
<GID>52</GID>
<name>IN_15</name></connection>
<connection>
<GID>53</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-76,20.5,-76</points>
<connection>
<GID>40</GID>
<name>IN_10</name></connection>
<connection>
<GID>2</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-51,20.5,-51</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1212 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-110,-62,-105</points>
<intersection>-110 1</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-110,-62,-110</points>
<connection>
<GID>1088</GID>
<name>OUT_1</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62,-105,-61,-105</points>
<connection>
<GID>1087</GID>
<name>IN_1</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>399 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-75,128.5,-75</points>
<connection>
<GID>55</GID>
<name>OUT_11</name></connection>
<connection>
<GID>54</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-50,20.5,-50</points>
<connection>
<GID>16</GID>
<name>IN_2</name></connection>
<connection>
<GID>10</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-74,20.5,-74</points>
<connection>
<GID>40</GID>
<name>IN_12</name></connection>
<connection>
<GID>2</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-44,117.5,-44</points>
<connection>
<GID>45</GID>
<name>OUT_8</name></connection>
<connection>
<GID>53</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>30 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-49,20.5,-49</points>
<connection>
<GID>16</GID>
<name>IN_3</name></connection>
<connection>
<GID>10</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>513 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>11,-153,11,-1</points>
<intersection>-153 32</intersection>
<intersection>-130 9</intersection>
<intersection>-89 10</intersection>
<intersection>-55 1</intersection>
<intersection>-1 25</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>5.5,-55,88,-55</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>11 0</intersection>
<intersection>24.5 13</intersection>
<intersection>88 27</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>11,-130,88,-130</points>
<intersection>11 0</intersection>
<intersection>24.5 17</intersection>
<intersection>88 33</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>11,-89,98.5,-89</points>
<intersection>11 0</intersection>
<intersection>24.5 15</intersection>
<intersection>98.5 14</intersection></hsegment>
<vsegment>
<ID>13</ID>
<points>24.5,-55,24.5,-54</points>
<connection>
<GID>10</GID>
<name>clock</name></connection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>14</ID>
<points>98.5,-89,98.5,-88</points>
<connection>
<GID>47</GID>
<name>clock</name></connection>
<intersection>-89 10</intersection></vsegment>
<vsegment>
<ID>15</ID>
<points>24.5,-89,24.5,-88</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>-89 10</intersection></vsegment>
<vsegment>
<ID>17</ID>
<points>24.5,-130,24.5,-129</points>
<connection>
<GID>29</GID>
<name>clock</name></connection>
<intersection>-130 9</intersection></vsegment>
<hsegment>
<ID>25</ID>
<points>11,-1,84,-1</points>
<intersection>11 0</intersection>
<intersection>84 28</intersection></hsegment>
<vsegment>
<ID>27</ID>
<points>88,-55,88,-54</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>-55 1</intersection></vsegment>
<vsegment>
<ID>28</ID>
<points>84,-10.5,84,-1</points>
<intersection>-10.5 29</intersection>
<intersection>-1 25</intersection></vsegment>
<hsegment>
<ID>29</ID>
<points>83,-10.5,84,-10.5</points>
<connection>
<GID>8</GID>
<name>write_clock</name></connection>
<intersection>84 28</intersection></hsegment>
<hsegment>
<ID>32</ID>
<points>11,-153,86.5,-153</points>
<intersection>11 0</intersection>
<intersection>86.5 39</intersection></hsegment>
<vsegment>
<ID>33</ID>
<points>88,-130,88,-129</points>
<connection>
<GID>13</GID>
<name>clock</name></connection>
<intersection>-130 9</intersection></vsegment>
<vsegment>
<ID>39</ID>
<points>86.5,-153,86.5,-152</points>
<connection>
<GID>116</GID>
<name>clock</name></connection>
<intersection>-153 32</intersection></vsegment></shape></wire>
<wire>
<ID>1208 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62,-100,-62,-95</points>
<intersection>-100 2</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-95,-62,-95</points>
<connection>
<GID>1086</GID>
<name>OUT_2</name></connection>
<intersection>-62 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62,-100,-61,-100</points>
<connection>
<GID>1087</GID>
<name>IN_6</name></connection>
<intersection>-62 0</intersection></hsegment></shape></wire>
<wire>
<ID>212 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-78,20.5,-78</points>
<connection>
<GID>40</GID>
<name>IN_8</name></connection>
<connection>
<GID>2</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>542 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-39,24.5,-34.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43,-52,43,-17.5</points>
<intersection>-52 2</intersection>
<intersection>-17.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-17.5,65,-17.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_0</name></connection>
<intersection>43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-52,54,-52</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>43 0</intersection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-51,42.5,-16.5</points>
<intersection>-51 2</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-16.5,65,-16.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_1</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-51,54,-51</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>10</GID>
<name>OUT_1</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38,-42,38,-7.5</points>
<intersection>-42 2</intersection>
<intersection>-7.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-7.5,65,-7.5</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_10</name></connection>
<intersection>38 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-42,54,-42</points>
<connection>
<GID>20</GID>
<name>IN_10</name></connection>
<connection>
<GID>10</GID>
<name>OUT_10</name></connection>
<intersection>38 0</intersection></hsegment></shape></wire>
<wire>
<ID>489 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-63,-46,-63</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37.5,-41,37.5,-6.5</points>
<intersection>-41 2</intersection>
<intersection>-6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-6.5,65,-6.5</points>
<connection>
<GID>82</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_11</name></connection>
<intersection>37.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-41,54,-41</points>
<connection>
<GID>20</GID>
<name>IN_11</name></connection>
<connection>
<GID>10</GID>
<name>OUT_11</name></connection>
<intersection>37.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42,-50,42,-15.5</points>
<intersection>-50 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-15.5,65,-15.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_2</name></connection>
<intersection>42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-50,54,-50</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<connection>
<GID>10</GID>
<name>OUT_2</name></connection>
<intersection>42 0</intersection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-49,41.5,-14.5</points>
<intersection>-49 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-14.5,65,-14.5</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_3</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-49,54,-49</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<connection>
<GID>10</GID>
<name>OUT_3</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41,-48,41,-13.5</points>
<intersection>-48 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-13.5,65,-13.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_4</name></connection>
<intersection>41 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-48,54,-48</points>
<connection>
<GID>20</GID>
<name>IN_4</name></connection>
<connection>
<GID>10</GID>
<name>OUT_4</name></connection>
<intersection>41 0</intersection></hsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-47,40.5,-12.5</points>
<intersection>-47 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-12.5,65,-12.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_5</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-47,54,-47</points>
<connection>
<GID>20</GID>
<name>IN_5</name></connection>
<connection>
<GID>10</GID>
<name>OUT_5</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40,-46,40,-11.5</points>
<intersection>-46 2</intersection>
<intersection>-11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-11.5,65,-11.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_6</name></connection>
<intersection>40 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-46,54,-46</points>
<connection>
<GID>20</GID>
<name>IN_6</name></connection>
<connection>
<GID>10</GID>
<name>OUT_6</name></connection>
<intersection>40 0</intersection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-45,39.5,-10.5</points>
<intersection>-45 2</intersection>
<intersection>-10.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-10.5,65,-10.5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_7</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-45,54,-45</points>
<connection>
<GID>20</GID>
<name>IN_7</name></connection>
<connection>
<GID>10</GID>
<name>OUT_7</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39,-44,39,-9.5</points>
<intersection>-44 2</intersection>
<intersection>-9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22.5,-9.5,65,-9.5</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_8</name></connection>
<intersection>39 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-44,54,-44</points>
<connection>
<GID>20</GID>
<name>IN_8</name></connection>
<connection>
<GID>10</GID>
<name>OUT_8</name></connection>
<intersection>39 0</intersection></hsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-43,38.5,-8.5</points>
<intersection>-43 2</intersection>
<intersection>-8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30.5,-8.5,65,-8.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>8</GID>
<name>ADDRESS_9</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>30.5,-43,54,-43</points>
<connection>
<GID>20</GID>
<name>IN_9</name></connection>
<connection>
<GID>10</GID>
<name>OUT_9</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1210 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-106,-63,-103</points>
<intersection>-106 1</intersection>
<intersection>-103 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-106,-63,-106</points>
<connection>
<GID>1088</GID>
<name>OUT_3</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-103,-61,-103</points>
<connection>
<GID>1087</GID>
<name>IN_3</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>214 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-86,20.5,-86</points>
<connection>
<GID>40</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-43,117.5,-43</points>
<connection>
<GID>45</GID>
<name>OUT_9</name></connection>
<connection>
<GID>53</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>557 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-76,54,-76</points>
<connection>
<GID>32</GID>
<name>IN_10</name></connection>
<connection>
<GID>2</GID>
<name>OUT_10</name></connection>
<intersection>34.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34.5,-101,34.5,-76</points>
<intersection>-101 4</intersection>
<intersection>-76 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34.5,-101,40,-101</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>34.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>219 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-85,20.5,-85</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>370 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-44,128.5,-44</points>
<connection>
<GID>52</GID>
<name>IN_8</name></connection>
<connection>
<GID>53</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>217 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-73,20.5,-73</points>
<connection>
<GID>40</GID>
<name>IN_13</name></connection>
<connection>
<GID>2</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>218 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-72,20.5,-72</points>
<connection>
<GID>40</GID>
<name>IN_14</name></connection>
<connection>
<GID>2</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>210 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-71,20.5,-71</points>
<connection>
<GID>40</GID>
<name>IN_15</name></connection>
<connection>
<GID>2</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>368 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-50,128.5,-50</points>
<connection>
<GID>52</GID>
<name>IN_2</name></connection>
<connection>
<GID>53</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>545 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-34,56,-34</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>56 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>56,-35.5,56,-34</points>
<connection>
<GID>20</GID>
<name>ENABLE_0</name></connection>
<intersection>-34 1</intersection></vsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-84,20.5,-84</points>
<connection>
<GID>40</GID>
<name>IN_2</name></connection>
<connection>
<GID>2</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>550 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-83,54,-83</points>
<connection>
<GID>32</GID>
<name>IN_3</name></connection>
<connection>
<GID>2</GID>
<name>OUT_3</name></connection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-94,38,-83</points>
<intersection>-94 4</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38,-94,48.5,-94</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>220 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-83,20.5,-83</points>
<connection>
<GID>40</GID>
<name>IN_3</name></connection>
<connection>
<GID>2</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1209 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,-99,-61.5,-93</points>
<intersection>-99 3</intersection>
<intersection>-93 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-93,-61.5,-93</points>
<connection>
<GID>1086</GID>
<name>OUT_3</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-61.5,-99,-61,-99</points>
<connection>
<GID>1087</GID>
<name>IN_7</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>366 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-47,128.5,-47</points>
<connection>
<GID>52</GID>
<name>IN_5</name></connection>
<connection>
<GID>53</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>213 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-82,20.5,-82</points>
<connection>
<GID>40</GID>
<name>IN_4</name></connection>
<connection>
<GID>2</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>215 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-81,20.5,-81</points>
<connection>
<GID>40</GID>
<name>IN_5</name></connection>
<connection>
<GID>2</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>554 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-79,54,-79</points>
<connection>
<GID>32</GID>
<name>IN_7</name></connection>
<connection>
<GID>2</GID>
<name>OUT_7</name></connection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-98,36,-79</points>
<intersection>-98 4</intersection>
<intersection>-79 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-98,48.5,-98</points>
<connection>
<GID>92</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-80,20.5,-80</points>
<connection>
<GID>40</GID>
<name>IN_6</name></connection>
<connection>
<GID>2</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>372 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-40,128.5,-40</points>
<connection>
<GID>52</GID>
<name>IN_12</name></connection>
<connection>
<GID>53</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>549 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-84,54,-84</points>
<connection>
<GID>32</GID>
<name>IN_2</name></connection>
<connection>
<GID>2</GID>
<name>OUT_2</name></connection>
<intersection>38.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38.5,-93,38.5,-84</points>
<intersection>-93 4</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>38.5,-93,40,-93</points>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>38.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>211 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-79,20.5,-79</points>
<connection>
<GID>40</GID>
<name>IN_7</name></connection>
<connection>
<GID>2</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>546 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-35.5,119.5,-34</points>
<connection>
<GID>53</GID>
<name>ENABLE_0</name></connection>
<intersection>-34 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>118,-34,119.5,-34</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>216 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-77,20.5,-77</points>
<connection>
<GID>40</GID>
<name>IN_9</name></connection>
<connection>
<GID>2</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>582 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-91,26.5,-88</points>
<connection>
<GID>2</GID>
<name>clear</name></connection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-91,26.5,-91</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>404 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-72,128.5,-72</points>
<connection>
<GID>55</GID>
<name>OUT_14</name></connection>
<connection>
<GID>54</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>581 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-69,25.5,-65</points>
<connection>
<GID>2</GID>
<name>count_enable</name></connection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>24.5,-65,25.5,-65</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>373 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-43,128.5,-43</points>
<connection>
<GID>52</GID>
<name>IN_9</name></connection>
<connection>
<GID>53</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>580 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-69,24.5,-67.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>398 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-78,128.5,-78</points>
<connection>
<GID>55</GID>
<name>OUT_8</name></connection>
<connection>
<GID>54</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>547 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-86,54,-86</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>39.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>39.5,-91,39.5,-86</points>
<intersection>-91 7</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>39.5,-91,40,-91</points>
<connection>
<GID>84</GID>
<name>IN_0</name></connection>
<intersection>39.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>548 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-85,54,-85</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>OUT_1</name></connection>
<intersection>39 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>39,-92,39,-85</points>
<intersection>-92 4</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>39,-92,48.5,-92</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<intersection>39 3</intersection></hsegment></shape></wire>
<wire>
<ID>228 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-116,20.5,-116</points>
<connection>
<GID>29</GID>
<name>IN_11</name></connection>
<connection>
<GID>41</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>558 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-75,54,-75</points>
<connection>
<GID>32</GID>
<name>IN_11</name></connection>
<connection>
<GID>2</GID>
<name>OUT_11</name></connection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-102,34,-75</points>
<intersection>-102 4</intersection>
<intersection>-75 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>34,-102,48.5,-102</points>
<connection>
<GID>96</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection></hsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-81,128.5,-81</points>
<connection>
<GID>55</GID>
<name>OUT_5</name></connection>
<connection>
<GID>54</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>559 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-74,54,-74</points>
<connection>
<GID>32</GID>
<name>IN_12</name></connection>
<connection>
<GID>2</GID>
<name>OUT_12</name></connection>
<intersection>33.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33.5,-103,33.5,-74</points>
<intersection>-103 4</intersection>
<intersection>-74 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33.5,-103,40,-103</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>33.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>560 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-73,54,-73</points>
<connection>
<GID>32</GID>
<name>IN_13</name></connection>
<connection>
<GID>2</GID>
<name>OUT_13</name></connection>
<intersection>33 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>33,-104,33,-73</points>
<intersection>-104 4</intersection>
<intersection>-73 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>33,-104,48.5,-104</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>33 3</intersection></hsegment></shape></wire>
<wire>
<ID>239 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-120,20.5,-120</points>
<connection>
<GID>29</GID>
<name>IN_7</name></connection>
<connection>
<GID>41</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>561 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-72,54,-72</points>
<connection>
<GID>32</GID>
<name>IN_14</name></connection>
<connection>
<GID>2</GID>
<name>OUT_14</name></connection>
<intersection>32.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32.5,-105,32.5,-72</points>
<intersection>-105 4</intersection>
<intersection>-72 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32.5,-105,40,-105</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>32.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>232 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-121,20.5,-121</points>
<connection>
<GID>29</GID>
<name>IN_6</name></connection>
<connection>
<GID>41</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>562 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-71,54,-71</points>
<connection>
<GID>32</GID>
<name>IN_15</name></connection>
<connection>
<GID>2</GID>
<name>OUT_15</name></connection>
<intersection>32 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>32,-106,32,-71</points>
<intersection>-106 4</intersection>
<intersection>-71 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>32,-106,48.5,-106</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>32 3</intersection></hsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-41,117.5,-41</points>
<connection>
<GID>45</GID>
<name>OUT_11</name></connection>
<connection>
<GID>53</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>551 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-82,54,-82</points>
<connection>
<GID>32</GID>
<name>IN_4</name></connection>
<connection>
<GID>2</GID>
<name>OUT_4</name></connection>
<intersection>37.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37.5,-95,37.5,-82</points>
<intersection>-95 4</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37.5,-95,40,-95</points>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>37.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>552 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-81,54,-81</points>
<connection>
<GID>32</GID>
<name>IN_5</name></connection>
<connection>
<GID>2</GID>
<name>OUT_5</name></connection>
<intersection>37 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>37,-96,37,-81</points>
<intersection>-96 4</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>37,-96,48.5,-96</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<intersection>37 3</intersection></hsegment></shape></wire>
<wire>
<ID>376 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-38,128.5,-38</points>
<connection>
<GID>52</GID>
<name>IN_14</name></connection>
<connection>
<GID>53</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>231 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-119,20.5,-119</points>
<connection>
<GID>29</GID>
<name>IN_8</name></connection>
<connection>
<GID>41</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>553 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-80,54,-80</points>
<connection>
<GID>32</GID>
<name>IN_6</name></connection>
<connection>
<GID>2</GID>
<name>OUT_6</name></connection>
<intersection>36.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-97,36.5,-80</points>
<intersection>-97 4</intersection>
<intersection>-80 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36.5,-97,40,-97</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>36.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>555 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-78,54,-78</points>
<connection>
<GID>32</GID>
<name>IN_8</name></connection>
<connection>
<GID>2</GID>
<name>OUT_8</name></connection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-99,35.5,-78</points>
<intersection>-99 4</intersection>
<intersection>-78 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35.5,-99,40,-99</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>35.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>907 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-52.5,-44.5,-51,-44.5</points>
<connection>
<GID>547</GID>
<name>OUT_0</name></connection>
<connection>
<GID>670</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>556 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>30.5,-77,54,-77</points>
<connection>
<GID>32</GID>
<name>IN_9</name></connection>
<connection>
<GID>2</GID>
<name>OUT_9</name></connection>
<intersection>35 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35,-100,35,-77</points>
<intersection>-100 4</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>35,-100,48.5,-100</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>35 3</intersection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-24,81.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-24,80.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_1</name></connection>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71.5,-24,71.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_10</name></connection>
<connection>
<GID>6</GID>
<name>IN_10</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_10</name></connection></vsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-24,70.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_11</name></connection>
<connection>
<GID>6</GID>
<name>IN_11</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_11</name></connection></vsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-24,69.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_12</name></connection>
<connection>
<GID>6</GID>
<name>IN_12</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_12</name></connection></vsegment></shape></wire>
<wire>
<ID>62 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68.5,-24,68.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_13</name></connection>
<connection>
<GID>6</GID>
<name>IN_13</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_13</name></connection></vsegment></shape></wire>
<wire>
<ID>72 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-24,67.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_14</name></connection>
<connection>
<GID>6</GID>
<name>IN_14</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_14</name></connection></vsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66.5,-24,66.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_15</name></connection>
<connection>
<GID>6</GID>
<name>IN_15</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_15</name></connection></vsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>79.5,-24,79.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_2</name></connection>
<connection>
<GID>6</GID>
<name>IN_2</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_2</name></connection></vsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78.5,-24,78.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_3</name></connection>
<connection>
<GID>6</GID>
<name>IN_3</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_3</name></connection></vsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>77.5,-24,77.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_4</name></connection>
<connection>
<GID>6</GID>
<name>IN_4</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_4</name></connection></vsegment></shape></wire>
<wire>
<ID>61 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>76.5,-24,76.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_5</name></connection>
<connection>
<GID>6</GID>
<name>IN_5</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_5</name></connection></vsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-24,75.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_6</name></connection>
<connection>
<GID>6</GID>
<name>IN_6</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_6</name></connection></vsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-24,74.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_7</name></connection>
<connection>
<GID>6</GID>
<name>IN_7</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_7</name></connection></vsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73.5,-24,73.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_8</name></connection>
<connection>
<GID>6</GID>
<name>IN_8</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_8</name></connection></vsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-24,72.5,-23</points>
<connection>
<GID>8</GID>
<name>DATA_OUT_9</name></connection>
<connection>
<GID>6</GID>
<name>IN_9</name></connection>
<connection>
<GID>8</GID>
<name>DATA_IN_9</name></connection></vsegment></shape></wire>
<wire>
<ID>708 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-13.5,84,-12.5</points>
<intersection>-13.5 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,-12.5,84,-12.5</points>
<connection>
<GID>8</GID>
<name>ENABLE_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>84,-13.5,85.5,-13.5</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>662 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-11.5,85.5,-11.5</points>
<connection>
<GID>8</GID>
<name>write_enable</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>307 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-52,84,-52</points>
<connection>
<GID>22</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>45</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-113,84,-113</points>
<connection>
<GID>17</GID>
<name>IN_14</name></connection>
<connection>
<GID>13</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>308 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-51,84,-51</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>45</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-126,117.5,-126</points>
<connection>
<GID>13</GID>
<name>OUT_1</name></connection>
<connection>
<GID>15</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>316 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-42,84,-42</points>
<connection>
<GID>22</GID>
<name>IN_10</name></connection>
<connection>
<GID>45</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>317 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-41,84,-41</points>
<connection>
<GID>22</GID>
<name>IN_11</name></connection>
<connection>
<GID>45</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-117,84,-117</points>
<connection>
<GID>17</GID>
<name>IN_10</name></connection>
<connection>
<GID>13</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>306 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-50,84,-50</points>
<connection>
<GID>22</GID>
<name>IN_2</name></connection>
<connection>
<GID>45</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>516 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-147,93,-147</points>
<connection>
<GID>116</GID>
<name>OUT_3</name></connection>
<connection>
<GID>139</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>309 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-49,84,-49</points>
<connection>
<GID>22</GID>
<name>IN_3</name></connection>
<connection>
<GID>45</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-124,117.5,-124</points>
<connection>
<GID>13</GID>
<name>OUT_3</name></connection>
<connection>
<GID>15</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>310 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-48,84,-48</points>
<connection>
<GID>22</GID>
<name>IN_4</name></connection>
<connection>
<GID>45</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>311 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-47,84,-47</points>
<connection>
<GID>22</GID>
<name>IN_5</name></connection>
<connection>
<GID>45</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-120,65,-120</points>
<connection>
<GID>35</GID>
<name>IN_7</name></connection>
<connection>
<GID>36</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>312 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-46,84,-46</points>
<connection>
<GID>22</GID>
<name>IN_6</name></connection>
<connection>
<GID>45</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>520 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-143,93,-143</points>
<connection>
<GID>116</GID>
<name>OUT_7</name></connection>
<connection>
<GID>139</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>313 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-45,84,-45</points>
<connection>
<GID>22</GID>
<name>IN_7</name></connection>
<connection>
<GID>45</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-120,117.5,-120</points>
<connection>
<GID>13</GID>
<name>OUT_7</name></connection>
<connection>
<GID>15</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>314 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-44,84,-44</points>
<connection>
<GID>22</GID>
<name>IN_8</name></connection>
<connection>
<GID>45</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>1216 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-102,-52,-102</points>
<connection>
<GID>1092</GID>
<name>IN_0</name></connection>
<connection>
<GID>1087</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>315 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,-43,84,-43</points>
<connection>
<GID>22</GID>
<name>IN_9</name></connection>
<connection>
<GID>45</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>237 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-127,20.5,-127</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>41</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-126,20.5,-126</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<connection>
<GID>41</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>570 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-79,117.5,-79</points>
<connection>
<GID>55</GID>
<name>IN_7</name></connection>
<connection>
<GID>47</GID>
<name>OUT_7</name></connection>
<intersection>110 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>110,-97.5,110,-79</points>
<intersection>-97.5 9</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>110,-97.5,123.5,-97.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>110 8</intersection></hsegment></shape></wire>
<wire>
<ID>240 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-117,20.5,-117</points>
<connection>
<GID>29</GID>
<name>IN_10</name></connection>
<connection>
<GID>41</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-51,117.5,-51</points>
<connection>
<GID>45</GID>
<name>OUT_1</name></connection>
<connection>
<GID>53</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>229 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-115,20.5,-115</points>
<connection>
<GID>29</GID>
<name>IN_12</name></connection>
<connection>
<GID>41</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>241 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-114,20.5,-114</points>
<connection>
<GID>29</GID>
<name>IN_13</name></connection>
<connection>
<GID>41</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>234 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-113,20.5,-113</points>
<connection>
<GID>29</GID>
<name>IN_14</name></connection>
<connection>
<GID>41</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>230 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-112,20.5,-112</points>
<connection>
<GID>29</GID>
<name>IN_15</name></connection>
<connection>
<GID>41</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>566 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-83,117.5,-83</points>
<connection>
<GID>55</GID>
<name>IN_3</name></connection>
<connection>
<GID>47</GID>
<name>OUT_3</name></connection>
<intersection>112 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>112,-93.5,112,-83</points>
<intersection>-93.5 6</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>112,-93.5,123.5,-93.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>112 5</intersection></hsegment></shape></wire>
<wire>
<ID>236 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-125,20.5,-125</points>
<connection>
<GID>29</GID>
<name>IN_2</name></connection>
<connection>
<GID>41</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>565 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-84,117.5,-84</points>
<connection>
<GID>55</GID>
<name>IN_2</name></connection>
<connection>
<GID>47</GID>
<name>OUT_2</name></connection>
<intersection>112.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>112.5,-92.5,112.5,-84</points>
<intersection>-92.5 9</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>112.5,-92.5,114,-92.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>112.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>227 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-124,20.5,-124</points>
<connection>
<GID>29</GID>
<name>IN_3</name></connection>
<connection>
<GID>41</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>573 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-76,117.5,-76</points>
<connection>
<GID>55</GID>
<name>IN_10</name></connection>
<connection>
<GID>47</GID>
<name>OUT_10</name></connection>
<intersection>108.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>108.5,-100.5,108.5,-76</points>
<intersection>-100.5 9</intersection>
<intersection>-76 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>108.5,-100.5,114,-100.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>108.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>235 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-123,20.5,-123</points>
<connection>
<GID>29</GID>
<name>IN_4</name></connection>
<connection>
<GID>41</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>238 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-122,20.5,-122</points>
<connection>
<GID>29</GID>
<name>IN_5</name></connection>
<connection>
<GID>41</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>233 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,-118,20.5,-118</points>
<connection>
<GID>29</GID>
<name>IN_9</name></connection>
<connection>
<GID>41</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>377 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-42,128.5,-42</points>
<connection>
<GID>52</GID>
<name>IN_10</name></connection>
<connection>
<GID>53</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>584 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24.5,-110,24.5,-108.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>971 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-76,94.5,-76</points>
<connection>
<GID>47</GID>
<name>IN_10</name></connection>
<connection>
<GID>861</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-127,54,-127</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>39.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>39.5,-132,39.5,-127</points>
<intersection>-132 11</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>39.5,-132,40,-132</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>39.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>968 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-86,94.5,-86</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<connection>
<GID>851</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-126,54,-126</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>OUT_1</name></connection>
<intersection>39 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>39,-133,39,-126</points>
<intersection>-133 11</intersection>
<intersection>-126 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>39,-133,48.5,-133</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>39 10</intersection></hsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-117,54,-117</points>
<connection>
<GID>36</GID>
<name>IN_10</name></connection>
<connection>
<GID>29</GID>
<name>OUT_10</name></connection>
<intersection>34.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>34.5,-142,34.5,-117</points>
<intersection>-142 11</intersection>
<intersection>-117 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>34.5,-142,40,-142</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>34.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>284 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-116,54,-116</points>
<connection>
<GID>36</GID>
<name>IN_11</name></connection>
<connection>
<GID>29</GID>
<name>OUT_11</name></connection>
<intersection>34 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>34,-143,34,-116</points>
<intersection>-143 11</intersection>
<intersection>-116 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>34,-143,48.5,-143</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>34 10</intersection></hsegment></shape></wire>
<wire>
<ID>133 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-115,128.5,-115</points>
<connection>
<GID>14</GID>
<name>IN_12</name></connection>
<connection>
<GID>15</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-115,54,-115</points>
<connection>
<GID>36</GID>
<name>IN_12</name></connection>
<connection>
<GID>29</GID>
<name>OUT_12</name></connection>
<intersection>33.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33.5,-144,33.5,-115</points>
<intersection>-144 11</intersection>
<intersection>-115 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>33.5,-144,40,-144</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>33.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-112,84,-112</points>
<connection>
<GID>17</GID>
<name>IN_15</name></connection>
<connection>
<GID>13</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-114,54,-114</points>
<connection>
<GID>36</GID>
<name>IN_13</name></connection>
<connection>
<GID>29</GID>
<name>OUT_13</name></connection>
<intersection>33 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>33,-145,33,-114</points>
<intersection>-145 11</intersection>
<intersection>-114 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>33,-145,48.5,-145</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<intersection>33 10</intersection></hsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-113,54,-113</points>
<connection>
<GID>36</GID>
<name>IN_14</name></connection>
<connection>
<GID>29</GID>
<name>OUT_14</name></connection>
<intersection>32.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>32.5,-146,32.5,-113</points>
<intersection>-146 11</intersection>
<intersection>-113 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>32.5,-146,40,-146</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>32.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>991 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-71,94.5,-71</points>
<connection>
<GID>47</GID>
<name>IN_15</name></connection>
<connection>
<GID>866</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-112,54,-112</points>
<connection>
<GID>36</GID>
<name>IN_15</name></connection>
<connection>
<GID>29</GID>
<name>OUT_15</name></connection>
<intersection>32 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>32,-147,32,-112</points>
<intersection>-147 11</intersection>
<intersection>-112 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>32,-147,48.5,-147</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>32 10</intersection></hsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-125,54,-125</points>
<connection>
<GID>36</GID>
<name>IN_2</name></connection>
<connection>
<GID>29</GID>
<name>OUT_2</name></connection>
<intersection>38.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>38.5,-134,38.5,-125</points>
<intersection>-134 11</intersection>
<intersection>-125 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>38.5,-134,40,-134</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>38.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-124,54,-124</points>
<connection>
<GID>36</GID>
<name>IN_3</name></connection>
<connection>
<GID>29</GID>
<name>OUT_3</name></connection>
<intersection>38 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>38,-135,38,-124</points>
<intersection>-135 11</intersection>
<intersection>-124 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>38,-135,48.5,-135</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>38 10</intersection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-123,54,-123</points>
<connection>
<GID>36</GID>
<name>IN_4</name></connection>
<connection>
<GID>29</GID>
<name>OUT_4</name></connection>
<intersection>37.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>37.5,-136,37.5,-123</points>
<intersection>-136 11</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>37.5,-136,40,-136</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>37.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>972 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-82,94.5,-82</points>
<connection>
<GID>47</GID>
<name>IN_4</name></connection>
<connection>
<GID>855</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-122,54,-122</points>
<connection>
<GID>36</GID>
<name>IN_5</name></connection>
<connection>
<GID>29</GID>
<name>OUT_5</name></connection>
<intersection>37 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>37,-137,37,-122</points>
<intersection>-137 11</intersection>
<intersection>-122 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>37,-137,48.5,-137</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>37 10</intersection></hsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-121,54,-121</points>
<connection>
<GID>36</GID>
<name>IN_6</name></connection>
<connection>
<GID>29</GID>
<name>OUT_6</name></connection>
<intersection>36.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>36.5,-138,36.5,-121</points>
<intersection>-138 11</intersection>
<intersection>-121 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>36.5,-138,40,-138</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>36.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-120,54,-120</points>
<connection>
<GID>36</GID>
<name>IN_7</name></connection>
<connection>
<GID>29</GID>
<name>OUT_7</name></connection>
<intersection>36 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>36,-139,36,-120</points>
<intersection>-139 11</intersection>
<intersection>-120 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>36,-139,48.5,-139</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>36 10</intersection></hsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-119,54,-119</points>
<connection>
<GID>36</GID>
<name>IN_8</name></connection>
<connection>
<GID>29</GID>
<name>OUT_8</name></connection>
<intersection>35.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>35.5,-140,35.5,-119</points>
<intersection>-140 11</intersection>
<intersection>-119 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>35.5,-140,40,-140</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>35.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-76,65,-76</points>
<connection>
<GID>32</GID>
<name>OUT_10</name></connection>
<connection>
<GID>31</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>30.5,-118,54,-118</points>
<connection>
<GID>36</GID>
<name>IN_9</name></connection>
<connection>
<GID>29</GID>
<name>OUT_9</name></connection>
<intersection>35 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>35,-141,35,-118</points>
<intersection>-141 11</intersection>
<intersection>-118 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>35,-141,48.5,-141</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>35 10</intersection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-86,65,-86</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<connection>
<GID>31</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>990 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-79,94.5,-79</points>
<connection>
<GID>47</GID>
<name>IN_7</name></connection>
<connection>
<GID>858</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-85,65,-85</points>
<connection>
<GID>32</GID>
<name>OUT_1</name></connection>
<connection>
<GID>31</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-75,65,-75</points>
<connection>
<GID>32</GID>
<name>OUT_11</name></connection>
<connection>
<GID>31</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>813 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-65.5,141.5,-65</points>
<connection>
<GID>304</GID>
<name>IN_4</name></connection>
<intersection>-65.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-65.5,143.5,-65.5</points>
<connection>
<GID>310</GID>
<name>IN_4</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-74,65,-74</points>
<connection>
<GID>32</GID>
<name>OUT_12</name></connection>
<connection>
<GID>31</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>986 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-77,94.5,-77</points>
<connection>
<GID>47</GID>
<name>IN_9</name></connection>
<connection>
<GID>860</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-73,65,-73</points>
<connection>
<GID>32</GID>
<name>OUT_13</name></connection>
<connection>
<GID>31</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-72,65,-72</points>
<connection>
<GID>32</GID>
<name>OUT_14</name></connection>
<connection>
<GID>31</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-71,65,-71</points>
<connection>
<GID>32</GID>
<name>OUT_15</name></connection>
<connection>
<GID>31</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>487 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-65.5,-51.5,-64</points>
<intersection>-65.5 5</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-64,-51,-64</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-54.5,-65.5,-51.5,-65.5</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-84,65,-84</points>
<connection>
<GID>32</GID>
<name>OUT_2</name></connection>
<connection>
<GID>31</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-83,65,-83</points>
<connection>
<GID>32</GID>
<name>OUT_3</name></connection>
<connection>
<GID>31</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-82,65,-82</points>
<connection>
<GID>32</GID>
<name>OUT_4</name></connection>
<connection>
<GID>31</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-81,65,-81</points>
<connection>
<GID>32</GID>
<name>OUT_5</name></connection>
<connection>
<GID>31</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-80,65,-80</points>
<connection>
<GID>32</GID>
<name>OUT_6</name></connection>
<connection>
<GID>31</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-79,65,-79</points>
<connection>
<GID>32</GID>
<name>OUT_7</name></connection>
<connection>
<GID>31</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-78,65,-78</points>
<connection>
<GID>32</GID>
<name>OUT_8</name></connection>
<connection>
<GID>31</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>844 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-59,141.5,-58.5</points>
<connection>
<GID>304</GID>
<name>IN_10</name></connection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-58.5,143.5,-58.5</points>
<connection>
<GID>312</GID>
<name>IN_2</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-77,65,-77</points>
<connection>
<GID>32</GID>
<name>OUT_9</name></connection>
<connection>
<GID>31</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>583 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-69.5,56,-68</points>
<connection>
<GID>32</GID>
<name>ENABLE_0</name></connection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-68,56,-68</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>486 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-51.5,-62,-51.5,-60.5</points>
<intersection>-62 1</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-51.5,-62,-51,-62</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>-51.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-52.5,-60.5,-51.5,-60.5</points>
<connection>
<GID>97</GID>
<name>CLK</name></connection>
<intersection>-51.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-127,65,-127</points>
<connection>
<GID>35</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-126,65,-126</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<connection>
<GID>36</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-117,65,-117</points>
<connection>
<GID>35</GID>
<name>IN_10</name></connection>
<connection>
<GID>36</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-116,65,-116</points>
<connection>
<GID>35</GID>
<name>IN_11</name></connection>
<connection>
<GID>36</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-115,65,-115</points>
<connection>
<GID>35</GID>
<name>IN_12</name></connection>
<connection>
<GID>36</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-114,65,-114</points>
<connection>
<GID>35</GID>
<name>IN_13</name></connection>
<connection>
<GID>36</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>865 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-57,141.5,-56.5</points>
<connection>
<GID>304</GID>
<name>IN_12</name></connection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-56.5,143.5,-56.5</points>
<connection>
<GID>312</GID>
<name>IN_4</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-113,65,-113</points>
<connection>
<GID>35</GID>
<name>IN_14</name></connection>
<connection>
<GID>36</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-112,65,-112</points>
<connection>
<GID>35</GID>
<name>IN_15</name></connection>
<connection>
<GID>36</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>1220 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-103,-43,-103</points>
<connection>
<GID>1087</GID>
<name>OUT_3</name></connection>
<connection>
<GID>1095</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-125,65,-125</points>
<connection>
<GID>35</GID>
<name>IN_2</name></connection>
<connection>
<GID>36</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-124,65,-124</points>
<connection>
<GID>35</GID>
<name>IN_3</name></connection>
<connection>
<GID>36</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-123,65,-123</points>
<connection>
<GID>35</GID>
<name>IN_4</name></connection>
<connection>
<GID>36</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-122,65,-122</points>
<connection>
<GID>35</GID>
<name>IN_5</name></connection>
<connection>
<GID>36</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1221 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-99,-43,-99</points>
<connection>
<GID>1097</GID>
<name>IN_0</name></connection>
<connection>
<GID>1087</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-121,65,-121</points>
<connection>
<GID>35</GID>
<name>IN_6</name></connection>
<connection>
<GID>36</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1222 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-101,-43,-101</points>
<connection>
<GID>1087</GID>
<name>OUT_5</name></connection>
<connection>
<GID>1096</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-119,65,-119</points>
<connection>
<GID>35</GID>
<name>IN_8</name></connection>
<connection>
<GID>36</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>58,-118,65,-118</points>
<connection>
<GID>35</GID>
<name>IN_9</name></connection>
<connection>
<GID>36</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-110,88,-108.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-109,56,-109</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>56 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>56,-110.5,56,-109</points>
<connection>
<GID>36</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>818 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-63.5,141.5,-63</points>
<connection>
<GID>304</GID>
<name>IN_6</name></connection>
<intersection>-63.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-63.5,143.5,-63.5</points>
<connection>
<GID>310</GID>
<name>IN_6</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>488 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-49,-60.5,-49,-59.5</points>
<connection>
<GID>101</GID>
<name>SEL_0</name></connection>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-110,89,-106</points>
<connection>
<GID>13</GID>
<name>count_enable</name></connection>
<intersection>-106 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-106,89,-106</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-115,117.5,-115</points>
<connection>
<GID>13</GID>
<name>OUT_12</name></connection>
<connection>
<GID>15</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>1219 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-105,-43,-105</points>
<connection>
<GID>1093</GID>
<name>IN_0</name></connection>
<connection>
<GID>1087</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>597 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-57,90,-54</points>
<connection>
<GID>45</GID>
<name>clear</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-57,90,-57</points>
<connection>
<GID>251</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>596 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,-39,89,-32</points>
<connection>
<GID>45</GID>
<name>count_enable</name></connection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-32,89,-32</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>595 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-39,88,-34.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<connection>
<GID>45</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-52,117.5,-52</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<connection>
<GID>53</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1206 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-63,-102,-63,-99</points>
<intersection>-102 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-99,-63,-99</points>
<connection>
<GID>1086</GID>
<name>OUT_0</name></connection>
<intersection>-63 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-63,-102,-61,-102</points>
<connection>
<GID>1087</GID>
<name>IN_4</name></connection>
<intersection>-63 0</intersection></hsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-42,117.5,-42</points>
<connection>
<GID>45</GID>
<name>OUT_10</name></connection>
<connection>
<GID>53</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-50,117.5,-50</points>
<connection>
<GID>45</GID>
<name>OUT_2</name></connection>
<connection>
<GID>53</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-47,117.5,-47</points>
<connection>
<GID>45</GID>
<name>OUT_5</name></connection>
<connection>
<GID>53</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>379 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-46,117.5,-46</points>
<connection>
<GID>45</GID>
<name>OUT_6</name></connection>
<connection>
<GID>53</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-45,117.5,-45</points>
<connection>
<GID>45</GID>
<name>OUT_7</name></connection>
<connection>
<GID>53</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>137 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-113,128.5,-113</points>
<connection>
<GID>14</GID>
<name>IN_14</name></connection>
<connection>
<GID>15</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>984 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-85,94.5,-85</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<connection>
<GID>852</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>987 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-75,94.5,-75</points>
<connection>
<GID>47</GID>
<name>IN_11</name></connection>
<connection>
<GID>862</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>973 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-74,94.5,-74</points>
<connection>
<GID>47</GID>
<name>IN_12</name></connection>
<connection>
<GID>863</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-116,84,-116</points>
<connection>
<GID>17</GID>
<name>IN_11</name></connection>
<connection>
<GID>13</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>988 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-73,94.5,-73</points>
<connection>
<GID>47</GID>
<name>IN_13</name></connection>
<connection>
<GID>864</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>975 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-72,94.5,-72</points>
<connection>
<GID>47</GID>
<name>IN_14</name></connection>
<connection>
<GID>865</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>969 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>93.5,-84,94.5,-84</points>
<connection>
<GID>47</GID>
<name>IN_2</name></connection>
<connection>
<GID>853</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>985 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-83,94.5,-83</points>
<connection>
<GID>47</GID>
<name>IN_3</name></connection>
<connection>
<GID>854</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>989 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>84.5,-81,94.5,-81</points>
<connection>
<GID>47</GID>
<name>IN_5</name></connection>
<connection>
<GID>856</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>593 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>100.5,-91,100.5,-88</points>
<connection>
<GID>47</GID>
<name>clear</name></connection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-91,100.5,-91</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>100.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>592 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>99.5,-69,99.5,-64.5</points>
<connection>
<GID>47</GID>
<name>count_enable</name></connection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>98.5,-64.5,99.5,-64.5</points>
<connection>
<GID>241</GID>
<name>IN_0</name></connection>
<intersection>99.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>591 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-69,98.5,-67.5</points>
<connection>
<GID>239</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>563 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-86,117.5,-86</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>OUT_0</name></connection>
<intersection>113.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>113.5,-90.5,113.5,-86</points>
<intersection>-90.5 12</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>113.5,-90.5,114,-90.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>113.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>564 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-85,117.5,-85</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<connection>
<GID>47</GID>
<name>OUT_1</name></connection>
<intersection>113 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>113,-91.5,113,-85</points>
<intersection>-91.5 9</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>113,-91.5,123.5,-91.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>113 8</intersection></hsegment></shape></wire>
<wire>
<ID>574 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-75,117.5,-75</points>
<connection>
<GID>55</GID>
<name>IN_11</name></connection>
<connection>
<GID>47</GID>
<name>OUT_11</name></connection>
<intersection>108 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>108,-101.5,108,-75</points>
<intersection>-101.5 9</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>108,-101.5,123.5,-101.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>108 8</intersection></hsegment></shape></wire>
<wire>
<ID>575 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-74,117.5,-74</points>
<connection>
<GID>55</GID>
<name>IN_12</name></connection>
<connection>
<GID>47</GID>
<name>OUT_12</name></connection>
<intersection>107.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>107.5,-102.5,107.5,-74</points>
<intersection>-102.5 13</intersection>
<intersection>-74 1</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>107.5,-102.5,114,-102.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>107.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>369 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-46,128.5,-46</points>
<connection>
<GID>52</GID>
<name>IN_6</name></connection>
<connection>
<GID>53</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>576 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-73,117.5,-73</points>
<connection>
<GID>55</GID>
<name>IN_13</name></connection>
<connection>
<GID>47</GID>
<name>OUT_13</name></connection>
<intersection>107 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>107,-103.5,107,-73</points>
<intersection>-103.5 9</intersection>
<intersection>-73 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>107,-103.5,123.5,-103.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>107 8</intersection></hsegment></shape></wire>
<wire>
<ID>400 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-74,128.5,-74</points>
<connection>
<GID>55</GID>
<name>OUT_12</name></connection>
<connection>
<GID>54</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>577 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-72,117.5,-72</points>
<connection>
<GID>55</GID>
<name>IN_14</name></connection>
<connection>
<GID>47</GID>
<name>OUT_14</name></connection>
<intersection>106.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>106.5,-104.5,106.5,-72</points>
<intersection>-104.5 9</intersection>
<intersection>-72 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>106.5,-104.5,114,-104.5</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>106.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>578 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-71,117.5,-71</points>
<connection>
<GID>55</GID>
<name>IN_15</name></connection>
<connection>
<GID>47</GID>
<name>OUT_15</name></connection>
<intersection>106 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>106,-105.5,106,-71</points>
<intersection>-105.5 9</intersection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>106,-105.5,123.5,-105.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>106 8</intersection></hsegment></shape></wire>
<wire>
<ID>402 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-71,128.5,-71</points>
<connection>
<GID>55</GID>
<name>OUT_15</name></connection>
<connection>
<GID>54</GID>
<name>IN_15</name></connection></hsegment></shape></wire>
<wire>
<ID>567 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-82,117.5,-82</points>
<connection>
<GID>55</GID>
<name>IN_4</name></connection>
<connection>
<GID>47</GID>
<name>OUT_4</name></connection>
<intersection>111.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>111.5,-94.5,111.5,-82</points>
<intersection>-94.5 9</intersection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>111.5,-94.5,114,-94.5</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>111.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>568 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-81,117.5,-81</points>
<connection>
<GID>55</GID>
<name>IN_5</name></connection>
<connection>
<GID>47</GID>
<name>OUT_5</name></connection>
<intersection>111 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>111,-95.5,111,-81</points>
<intersection>-95.5 9</intersection>
<intersection>-81 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>111,-95.5,123.5,-95.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>111 8</intersection></hsegment></shape></wire>
<wire>
<ID>569 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-80,117.5,-80</points>
<connection>
<GID>55</GID>
<name>IN_6</name></connection>
<connection>
<GID>47</GID>
<name>OUT_6</name></connection>
<intersection>110.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>110.5,-96.5,110.5,-80</points>
<intersection>-96.5 14</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>110.5,-96.5,114,-96.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>110.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>571 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-78,117.5,-78</points>
<connection>
<GID>55</GID>
<name>IN_8</name></connection>
<connection>
<GID>47</GID>
<name>OUT_8</name></connection>
<intersection>109.5 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>109.5,-98.5,109.5,-78</points>
<intersection>-98.5 9</intersection>
<intersection>-78 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>109.5,-98.5,114,-98.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>109.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>572 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,-77,117.5,-77</points>
<connection>
<GID>55</GID>
<name>IN_9</name></connection>
<connection>
<GID>47</GID>
<name>OUT_9</name></connection>
<intersection>109 8</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>109,-99.5,109,-77</points>
<intersection>-99.5 9</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>109,-99.5,123.5,-99.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>109 8</intersection></hsegment></shape></wire>
<wire>
<ID>1207 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-62.5,-101,-62.5,-97</points>
<intersection>-101 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-97,-62.5,-97</points>
<connection>
<GID>1086</GID>
<name>OUT_1</name></connection>
<intersection>-62.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62.5,-101,-61,-101</points>
<connection>
<GID>1087</GID>
<name>IN_5</name></connection>
<intersection>-62.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-150,83.5,-150</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-149,83.5,-149</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>521 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-146,93,-146</points>
<connection>
<GID>116</GID>
<name>OUT_4</name></connection>
<connection>
<GID>139</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-148,83.5,-148</points>
<connection>
<GID>116</GID>
<name>IN_2</name></connection>
<connection>
<GID>28</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-147,83.5,-147</points>
<connection>
<GID>116</GID>
<name>IN_3</name></connection>
<connection>
<GID>28</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-146,83.5,-146</points>
<connection>
<GID>116</GID>
<name>IN_4</name></connection>
<connection>
<GID>28</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-145,83.5,-145</points>
<connection>
<GID>116</GID>
<name>IN_5</name></connection>
<connection>
<GID>28</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-144,83.5,-144</points>
<connection>
<GID>116</GID>
<name>IN_6</name></connection>
<connection>
<GID>28</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82.5,-143,83.5,-143</points>
<connection>
<GID>116</GID>
<name>IN_7</name></connection>
<connection>
<GID>28</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>86.5,-141,86.5,-138.5</points>
<connection>
<GID>116</GID>
<name>load</name></connection>
<intersection>-138.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>86.5,-138.5,87.5,-138.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>86.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>514 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-150,93,-150</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<connection>
<GID>139</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>518 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-149,93,-149</points>
<connection>
<GID>116</GID>
<name>OUT_1</name></connection>
<connection>
<GID>139</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>515 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-148,93,-148</points>
<connection>
<GID>116</GID>
<name>OUT_2</name></connection>
<connection>
<GID>139</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>519 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-145,93,-145</points>
<connection>
<GID>116</GID>
<name>OUT_5</name></connection>
<connection>
<GID>139</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>517 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,-144,93,-144</points>
<connection>
<GID>116</GID>
<name>OUT_6</name></connection>
<connection>
<GID>139</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-52,128.5,-52</points>
<connection>
<GID>52</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-51,128.5,-51</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<connection>
<GID>53</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>371 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-41,128.5,-41</points>
<connection>
<GID>52</GID>
<name>IN_11</name></connection>
<connection>
<GID>53</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>375 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-39,128.5,-39</points>
<connection>
<GID>52</GID>
<name>IN_13</name></connection>
<connection>
<GID>53</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>1215 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-106,-52,-106</points>
<connection>
<GID>1094</GID>
<name>IN_0</name></connection>
<connection>
<GID>1087</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>364 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-49,128.5,-49</points>
<connection>
<GID>52</GID>
<name>IN_3</name></connection>
<connection>
<GID>53</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>365 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-48,128.5,-48</points>
<connection>
<GID>52</GID>
<name>IN_4</name></connection>
<connection>
<GID>53</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>367 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-45,128.5,-45</points>
<connection>
<GID>52</GID>
<name>IN_7</name></connection>
<connection>
<GID>53</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>594 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-69.5,119.5,-68</points>
<connection>
<GID>55</GID>
<name>ENABLE_0</name></connection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-68,119.5,-68</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-86,128.5,-86</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<connection>
<GID>54</GID>
<name>Bus_in_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1204 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-55.5,-74.5,-54.5,-74.5</points>
<connection>
<GID>1079</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1081</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-85,128.5,-85</points>
<connection>
<GID>55</GID>
<name>OUT_1</name></connection>
<connection>
<GID>54</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-84,128.5,-84</points>
<connection>
<GID>55</GID>
<name>OUT_2</name></connection>
<connection>
<GID>54</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-83,128.5,-83</points>
<connection>
<GID>55</GID>
<name>OUT_3</name></connection>
<connection>
<GID>54</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>843 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-61,141.5,-60.5</points>
<connection>
<GID>304</GID>
<name>IN_8</name></connection>
<intersection>-60.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-60.5,143.5,-60.5</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>864 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-60,141.5,-59.5</points>
<connection>
<GID>304</GID>
<name>IN_9</name></connection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-59.5,143.5,-59.5</points>
<connection>
<GID>312</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>863 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-58,141.5,-57.5</points>
<connection>
<GID>304</GID>
<name>IN_11</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-57.5,143.5,-57.5</points>
<connection>
<GID>312</GID>
<name>IN_3</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>839 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-56,141.5,-55.5</points>
<connection>
<GID>304</GID>
<name>IN_13</name></connection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-55.5,143.5,-55.5</points>
<connection>
<GID>312</GID>
<name>IN_5</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-117,117.5,-117</points>
<connection>
<GID>13</GID>
<name>OUT_10</name></connection>
<connection>
<GID>15</GID>
<name>IN_10</name></connection></hsegment></shape></wire>
<wire>
<ID>869 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-55,141.5,-54.5</points>
<connection>
<GID>304</GID>
<name>IN_14</name></connection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-54.5,143.5,-54.5</points>
<connection>
<GID>312</GID>
<name>IN_6</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>870 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-54,141.5,-53.5</points>
<connection>
<GID>304</GID>
<name>IN_15</name></connection>
<intersection>-53.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-53.5,143.5,-53.5</points>
<connection>
<GID>312</GID>
<name>IN_7</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-132,90,-129</points>
<connection>
<GID>13</GID>
<name>clear</name></connection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-132,90,-132</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>811 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-69.5,141.5,-69</points>
<connection>
<GID>304</GID>
<name>Bus_in_0</name></connection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-69.5,143.5,-69.5</points>
<connection>
<GID>310</GID>
<name>IN_0</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-127,84,-127</points>
<connection>
<GID>17</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-126,84,-126</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<connection>
<GID>13</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-115,84,-115</points>
<connection>
<GID>17</GID>
<name>IN_12</name></connection>
<connection>
<GID>13</GID>
<name>IN_12</name></connection></hsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-114,84,-114</points>
<connection>
<GID>17</GID>
<name>IN_13</name></connection>
<connection>
<GID>13</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-125,84,-125</points>
<connection>
<GID>17</GID>
<name>IN_2</name></connection>
<connection>
<GID>13</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-124,84,-124</points>
<connection>
<GID>17</GID>
<name>IN_3</name></connection>
<connection>
<GID>13</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>837 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-68.5,141.5,-68</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-68.5,143.5,-68.5</points>
<connection>
<GID>310</GID>
<name>IN_1</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-123,84,-123</points>
<connection>
<GID>17</GID>
<name>IN_4</name></connection>
<connection>
<GID>13</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-122,84,-122</points>
<connection>
<GID>17</GID>
<name>IN_5</name></connection>
<connection>
<GID>13</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-121,84,-121</points>
<connection>
<GID>17</GID>
<name>IN_6</name></connection>
<connection>
<GID>13</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-120,84,-120</points>
<connection>
<GID>17</GID>
<name>IN_7</name></connection>
<connection>
<GID>13</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-119,84,-119</points>
<connection>
<GID>17</GID>
<name>IN_8</name></connection>
<connection>
<GID>13</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>83,-118,84,-118</points>
<connection>
<GID>17</GID>
<name>IN_9</name></connection>
<connection>
<GID>13</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-127,117.5,-127</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-116,117.5,-116</points>
<connection>
<GID>13</GID>
<name>OUT_11</name></connection>
<connection>
<GID>15</GID>
<name>IN_11</name></connection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-114,117.5,-114</points>
<connection>
<GID>13</GID>
<name>OUT_13</name></connection>
<connection>
<GID>15</GID>
<name>IN_13</name></connection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-113,117.5,-113</points>
<connection>
<GID>13</GID>
<name>OUT_14</name></connection>
<connection>
<GID>15</GID>
<name>IN_14</name></connection></hsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-112,117.5,-112</points>
<connection>
<GID>15</GID>
<name>IN_15</name></connection>
<connection>
<GID>13</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-125,117.5,-125</points>
<connection>
<GID>13</GID>
<name>OUT_2</name></connection>
<connection>
<GID>15</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-123,117.5,-123</points>
<connection>
<GID>13</GID>
<name>OUT_4</name></connection>
<connection>
<GID>15</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-122,117.5,-122</points>
<connection>
<GID>13</GID>
<name>OUT_5</name></connection>
<connection>
<GID>15</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-121,117.5,-121</points>
<connection>
<GID>13</GID>
<name>OUT_6</name></connection>
<connection>
<GID>15</GID>
<name>IN_6</name></connection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-119,117.5,-119</points>
<connection>
<GID>13</GID>
<name>OUT_8</name></connection>
<connection>
<GID>15</GID>
<name>IN_8</name></connection></hsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94,-118,117.5,-118</points>
<connection>
<GID>13</GID>
<name>OUT_9</name></connection>
<connection>
<GID>15</GID>
<name>IN_9</name></connection></hsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-127,128.5,-127</points>
<connection>
<GID>14</GID>
<name>Bus_in_0</name></connection>
<connection>
<GID>15</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-126,128.5,-126</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>15</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>138 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-117,128.5,-117</points>
<connection>
<GID>14</GID>
<name>IN_10</name></connection>
<connection>
<GID>15</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>132 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-116,128.5,-116</points>
<connection>
<GID>14</GID>
<name>IN_11</name></connection>
<connection>
<GID>15</GID>
<name>OUT_11</name></connection></hsegment></shape></wire>
<wire>
<ID>136 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-114,128.5,-114</points>
<connection>
<GID>14</GID>
<name>IN_13</name></connection>
<connection>
<GID>15</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121.5,-112,128.5,-112</points>
<connection>
<GID>14</GID>
<name>IN_15</name></connection>
<connection>
<GID>15</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-125,128.5,-125</points>
<connection>
<GID>14</GID>
<name>IN_2</name></connection>
<connection>
<GID>15</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-124,128.5,-124</points>
<connection>
<GID>14</GID>
<name>IN_3</name></connection>
<connection>
<GID>15</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-123,128.5,-123</points>
<connection>
<GID>14</GID>
<name>IN_4</name></connection>
<connection>
<GID>15</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-122,128.5,-122</points>
<connection>
<GID>14</GID>
<name>IN_5</name></connection>
<connection>
<GID>15</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-121,128.5,-121</points>
<connection>
<GID>14</GID>
<name>IN_6</name></connection>
<connection>
<GID>15</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-120,128.5,-120</points>
<connection>
<GID>14</GID>
<name>IN_7</name></connection>
<connection>
<GID>15</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-119,128.5,-119</points>
<connection>
<GID>14</GID>
<name>IN_8</name></connection>
<connection>
<GID>15</GID>
<name>OUT_8</name></connection></hsegment></shape></wire>
<wire>
<ID>134 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>121.5,-118,128.5,-118</points>
<connection>
<GID>14</GID>
<name>IN_9</name></connection>
<connection>
<GID>15</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>119.5,-110.5,119.5,-109</points>
<connection>
<GID>15</GID>
<name>ENABLE_0</name></connection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-109,119.5,-109</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>119.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1223 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-58,-97,-58,-96</points>
<connection>
<GID>1098</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1087</GID>
<name>load</name></connection></vsegment></shape></wire>
<wire>
<ID>1218 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-104,-52,-104</points>
<connection>
<GID>1087</GID>
<name>OUT_2</name></connection>
<connection>
<GID>1089</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1217 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-53,-100,-52,-100</points>
<connection>
<GID>1087</GID>
<name>OUT_6</name></connection>
<connection>
<GID>1090</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1205 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-55.5,-78.5,-54.5,-78.5</points>
<connection>
<GID>1083</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1082</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>817 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-67.5,141.5,-67</points>
<connection>
<GID>304</GID>
<name>IN_2</name></connection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-67.5,143.5,-67.5</points>
<connection>
<GID>310</GID>
<name>IN_2</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>838 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-66.5,141.5,-66</points>
<connection>
<GID>304</GID>
<name>IN_3</name></connection>
<intersection>-66.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-66.5,143.5,-66.5</points>
<connection>
<GID>310</GID>
<name>IN_3</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>792 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-64.5,141.5,-64</points>
<connection>
<GID>304</GID>
<name>IN_5</name></connection>
<intersection>-64.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-64.5,143.5,-64.5</points>
<connection>
<GID>310</GID>
<name>IN_5</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>812 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>141.5,-62.5,141.5,-62</points>
<connection>
<GID>304</GID>
<name>IN_7</name></connection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>141.5,-62.5,143.5,-62.5</points>
<connection>
<GID>310</GID>
<name>IN_7</name></connection>
<intersection>141.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-131.975,-86.625,162.3,-235.25</PageViewport>
<gate>
<ID>197</ID>
<type>DA_FROM</type>
<position>-108,-127</position>
<input>
<ID>IN_0</ID>266 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR8</lparam></gate>
<gate>
<ID>177</ID>
<type>DE_TO</type>
<position>-84.5,-114.5</position>
<input>
<ID>IN_0</ID>251 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add5</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_AND2</type>
<position>74,-89</position>
<input>
<ID>IN_0</ID>447 </input>
<input>
<ID>IN_1</ID>446 </input>
<output>
<ID>OUT</ID>445 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>-108,-144</position>
<input>
<ID>IN_0</ID>263 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR12</lparam></gate>
<gate>
<ID>711</ID>
<type>DA_FROM</type>
<position>-42,-212</position>
<input>
<ID>IN_0</ID>851 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>190</ID>
<type>DA_FROM</type>
<position>-116,-94</position>
<input>
<ID>IN_0</ID>267 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR1</lparam></gate>
<gate>
<ID>198</ID>
<type>DA_FROM</type>
<position>-116,-128</position>
<input>
<ID>IN_0</ID>271 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR9</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>-116,-111</position>
<input>
<ID>IN_0</ID>273 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR5</lparam></gate>
<gate>
<ID>465</ID>
<type>DA_FROM</type>
<position>-3,-128.5</position>
<input>
<ID>IN_0</ID>614 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR5</lparam></gate>
<gate>
<ID>218</ID>
<type>DA_FROM</type>
<position>-117.5,-137</position>
<input>
<ID>IN_0</ID>318 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo11</lparam></gate>
<gate>
<ID>154</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-101,-98</position>
<input>
<ID>IN_0</ID>293 </input>
<input>
<ID>IN_1</ID>301 </input>
<input>
<ID>IN_2</ID>294 </input>
<input>
<ID>IN_3</ID>302 </input>
<input>
<ID>IN_B_0</ID>261 </input>
<input>
<ID>IN_B_1</ID>267 </input>
<input>
<ID>IN_B_2</ID>262 </input>
<input>
<ID>IN_B_3</ID>268 </input>
<output>
<ID>OUT_0</ID>245 </output>
<output>
<ID>OUT_1</ID>254 </output>
<output>
<ID>OUT_2</ID>246 </output>
<output>
<ID>OUT_3</ID>253 </output>
<input>
<ID>carry_in</ID>209 </input>
<output>
<ID>carry_out</ID>206 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>449</ID>
<type>DA_FROM</type>
<position>68,-147.5</position>
<input>
<ID>IN_0</ID>600 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>522</ID>
<type>AA_AND2</type>
<position>74,-183.5</position>
<input>
<ID>IN_0</ID>728 </input>
<input>
<ID>IN_1</ID>727 </input>
<output>
<ID>OUT</ID>726 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>-116,-96</position>
<input>
<ID>IN_0</ID>268 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR3</lparam></gate>
<gate>
<ID>526</ID>
<type>DA_FROM</type>
<position>68,-182.5</position>
<input>
<ID>IN_0</ID>728 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>196</ID>
<type>DA_FROM</type>
<position>-116,-113</position>
<input>
<ID>IN_0</ID>290 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR7</lparam></gate>
<gate>
<ID>530</ID>
<type>AA_AND2</type>
<position>-36,-168.5</position>
<input>
<ID>IN_0</ID>665 </input>
<input>
<ID>IN_1</ID>664 </input>
<output>
<ID>OUT</ID>663 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>DA_FROM</type>
<position>-116,-130</position>
<input>
<ID>IN_0</ID>272 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR11</lparam></gate>
<gate>
<ID>534</ID>
<type>DA_FROM</type>
<position>-58,-170.5</position>
<input>
<ID>IN_0</ID>667 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo8</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>-116,-147</position>
<input>
<ID>IN_0</ID>270 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR15</lparam></gate>
<gate>
<ID>316</ID>
<type>FF_GND</type>
<position>-27.5,-100</position>
<output>
<ID>OUT_0</ID>414 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>155</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-101,-115</position>
<input>
<ID>IN_0</ID>291 </input>
<input>
<ID>IN_1</ID>300 </input>
<input>
<ID>IN_2</ID>292 </input>
<input>
<ID>IN_3</ID>299 </input>
<input>
<ID>IN_B_0</ID>259 </input>
<input>
<ID>IN_B_1</ID>273 </input>
<input>
<ID>IN_B_2</ID>260 </input>
<input>
<ID>IN_B_3</ID>290 </input>
<output>
<ID>OUT_0</ID>244 </output>
<output>
<ID>OUT_1</ID>251 </output>
<output>
<ID>OUT_2</ID>243 </output>
<output>
<ID>OUT_3</ID>252 </output>
<input>
<ID>carry_in</ID>206 </input>
<output>
<ID>carry_out</ID>207 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>550</ID>
<type>DA_FROM</type>
<position>-42,-189.5</position>
<input>
<ID>IN_0</ID>685 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo9</lparam></gate>
<gate>
<ID>220</ID>
<type>DA_FROM</type>
<position>-108,-151</position>
<input>
<ID>IN_0</ID>296 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo12</lparam></gate>
<gate>
<ID>156</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-101,-132</position>
<input>
<ID>IN_0</ID>298 </input>
<input>
<ID>IN_1</ID>305 </input>
<input>
<ID>IN_2</ID>297 </input>
<input>
<ID>IN_3</ID>318 </input>
<input>
<ID>IN_B_0</ID>266 </input>
<input>
<ID>IN_B_1</ID>271 </input>
<input>
<ID>IN_B_2</ID>265 </input>
<input>
<ID>IN_B_3</ID>272 </input>
<output>
<ID>OUT_0</ID>247 </output>
<output>
<ID>OUT_1</ID>256 </output>
<output>
<ID>OUT_2</ID>248 </output>
<output>
<ID>OUT_3</ID>257 </output>
<input>
<ID>carry_in</ID>207 </input>
<output>
<ID>carry_out</ID>208 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>157</ID>
<type>AE_FULLADDER_4BIT</type>
<position>-101,-149</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>304 </input>
<input>
<ID>IN_2</ID>295 </input>
<input>
<ID>IN_3</ID>303 </input>
<input>
<ID>IN_B_0</ID>263 </input>
<input>
<ID>IN_B_1</ID>269 </input>
<input>
<ID>IN_B_2</ID>264 </input>
<input>
<ID>IN_B_3</ID>270 </input>
<output>
<ID>OUT_0</ID>249 </output>
<output>
<ID>OUT_1</ID>258 </output>
<output>
<ID>OUT_2</ID>250 </output>
<output>
<ID>OUT_3</ID>255 </output>
<input>
<ID>carry_in</ID>208 </input>
<output>
<ID>carry_out</ID>348 </output>
<gparam>angle 90</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>159</ID>
<type>FF_GND</type>
<position>-100.5,-89</position>
<output>
<ID>OUT_0</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>-94,-96.5</position>
<input>
<ID>IN_0</ID>245 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add0</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>-84.5,-97.5</position>
<input>
<ID>IN_0</ID>254 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add1</lparam></gate>
<gate>
<ID>164</ID>
<type>DE_TO</type>
<position>-94,-98.5</position>
<input>
<ID>IN_0</ID>246 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add2</lparam></gate>
<gate>
<ID>166</ID>
<type>DE_TO</type>
<position>-84.5,-99.5</position>
<input>
<ID>IN_0</ID>253 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add3</lparam></gate>
<gate>
<ID>176</ID>
<type>DE_TO</type>
<position>-94,-113.5</position>
<input>
<ID>IN_0</ID>244 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add4</lparam></gate>
<gate>
<ID>178</ID>
<type>DE_TO</type>
<position>-94,-115.5</position>
<input>
<ID>IN_0</ID>243 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add6</lparam></gate>
<gate>
<ID>179</ID>
<type>DE_TO</type>
<position>-84.5,-116.5</position>
<input>
<ID>IN_0</ID>252 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add7</lparam></gate>
<gate>
<ID>1048</ID>
<type>DE_TO</type>
<position>-95,-161</position>
<input>
<ID>IN_0</ID>1177 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Cout</lparam></gate>
<gate>
<ID>180</ID>
<type>DE_TO</type>
<position>-94,-130.5</position>
<input>
<ID>IN_0</ID>247 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add8</lparam></gate>
<gate>
<ID>181</ID>
<type>DE_TO</type>
<position>-84.5,-131.5</position>
<input>
<ID>IN_0</ID>256 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add9</lparam></gate>
<gate>
<ID>182</ID>
<type>DE_TO</type>
<position>-94,-132.5</position>
<input>
<ID>IN_0</ID>248 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add10</lparam></gate>
<gate>
<ID>183</ID>
<type>DE_TO</type>
<position>-84.5,-133.5</position>
<input>
<ID>IN_0</ID>257 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add11</lparam></gate>
<gate>
<ID>184</ID>
<type>DE_TO</type>
<position>-94,-147.5</position>
<input>
<ID>IN_0</ID>249 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add12</lparam></gate>
<gate>
<ID>185</ID>
<type>DE_TO</type>
<position>-84.5,-148.5</position>
<input>
<ID>IN_0</ID>258 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add13</lparam></gate>
<gate>
<ID>186</ID>
<type>DE_TO</type>
<position>-94,-149.5</position>
<input>
<ID>IN_0</ID>250 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add14</lparam></gate>
<gate>
<ID>187</ID>
<type>DE_TO</type>
<position>-84.5,-150.5</position>
<input>
<ID>IN_0</ID>255 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add15</lparam></gate>
<gate>
<ID>189</ID>
<type>DA_FROM</type>
<position>-108,-93</position>
<input>
<ID>IN_0</ID>261 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR0</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>-108,-95</position>
<input>
<ID>IN_0</ID>262 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR2</lparam></gate>
<gate>
<ID>346</ID>
<type>DA_FROM</type>
<position>13,-120</position>
<input>
<ID>IN_0</ID>439 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR1</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>-108,-110</position>
<input>
<ID>IN_0</ID>259 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR4</lparam></gate>
<gate>
<ID>533</ID>
<type>DA_FROM</type>
<position>-58,-168.5</position>
<input>
<ID>IN_0</ID>666 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR8</lparam></gate>
<gate>
<ID>356</ID>
<type>DA_FROM</type>
<position>68,-88</position>
<input>
<ID>IN_0</ID>447 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>195</ID>
<type>DA_FROM</type>
<position>-108,-112</position>
<input>
<ID>IN_0</ID>260 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR6</lparam></gate>
<gate>
<ID>344</ID>
<type>DA_FROM</type>
<position>13,-118</position>
<input>
<ID>IN_0</ID>437 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>199</ID>
<type>DA_FROM</type>
<position>-108,-129</position>
<input>
<ID>IN_0</ID>265 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR10</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>-116,-145</position>
<input>
<ID>IN_0</ID>269 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR13</lparam></gate>
<gate>
<ID>541</ID>
<type>AE_SMALL_INVERTER</type>
<position>-51,-184.5</position>
<input>
<ID>IN_0</ID>667 </input>
<output>
<ID>OUT_0</ID>675 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>364</ID>
<type>AA_AND2</type>
<position>74,-104</position>
<input>
<ID>IN_0</ID>458 </input>
<input>
<ID>IN_1</ID>457 </input>
<output>
<ID>OUT</ID>456 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>-108,-146</position>
<input>
<ID>IN_0</ID>264 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR14</lparam></gate>
<gate>
<ID>206</ID>
<type>DA_FROM</type>
<position>-108,-100</position>
<input>
<ID>IN_0</ID>293 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>529</ID>
<type>DE_OR8</type>
<position>-23.5,-183.5</position>
<input>
<ID>IN_0</ID>684 </input>
<input>
<ID>IN_1</ID>663 </input>
<input>
<ID>IN_2</ID>671 </input>
<input>
<ID>IN_3</ID>672 </input>
<input>
<ID>IN_4</ID>871 </input>
<input>
<ID>IN_5</ID>679 </input>
<input>
<ID>IN_6</ID>677 </input>
<input>
<ID>IN_7</ID>674 </input>
<output>
<ID>OUT</ID>668 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>352</ID>
<type>DE_TO</type>
<position>93.5,-104</position>
<input>
<ID>IN_0</ID>450 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi2</lparam></gate>
<gate>
<ID>207</ID>
<type>DA_FROM</type>
<position>-117.5,-101</position>
<input>
<ID>IN_0</ID>301 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo1</lparam></gate>
<gate>
<ID>538</ID>
<type>AA_AND2</type>
<position>-36,-178.5</position>
<input>
<ID>IN_0</ID>673 </input>
<input>
<ID>IN_1</ID>666 </input>
<output>
<ID>OUT</ID>672 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>DA_FROM</type>
<position>-108,-102</position>
<input>
<ID>IN_0</ID>294 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo2</lparam></gate>
<gate>
<ID>362</ID>
<type>AA_AND2</type>
<position>74,-99</position>
<input>
<ID>IN_0</ID>455 </input>
<input>
<ID>IN_1</ID>448 </input>
<output>
<ID>OUT</ID>454 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>DA_FROM</type>
<position>-117.5,-103</position>
<input>
<ID>IN_0</ID>302 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo3</lparam></gate>
<gate>
<ID>210</ID>
<type>DA_FROM</type>
<position>-108,-117</position>
<input>
<ID>IN_0</ID>291 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo4</lparam></gate>
<gate>
<ID>372</ID>
<type>AA_AND2</type>
<position>74,-119</position>
<input>
<ID>IN_0</ID>463 </input>
<input>
<ID>IN_1</ID>465 </input>
<output>
<ID>OUT</ID>464 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>DA_FROM</type>
<position>-117.5,-118</position>
<input>
<ID>IN_0</ID>300 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo5</lparam></gate>
<gate>
<ID>542</ID>
<type>DA_FROM</type>
<position>-42,-182.5</position>
<input>
<ID>IN_0</ID>676 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>212</ID>
<type>DA_FROM</type>
<position>-108,-119</position>
<input>
<ID>IN_0</ID>292 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo6</lparam></gate>
<gate>
<ID>366</ID>
<type>DA_FROM</type>
<position>68,-103</position>
<input>
<ID>IN_0</ID>458 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>213</ID>
<type>DA_FROM</type>
<position>-117.5,-120</position>
<input>
<ID>IN_0</ID>299 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo7</lparam></gate>
<gate>
<ID>214</ID>
<type>DA_FROM</type>
<position>-108,-134</position>
<input>
<ID>IN_0</ID>298 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo8</lparam></gate>
<gate>
<ID>537</ID>
<type>DA_FROM</type>
<position>-42,-174.5</position>
<input>
<ID>IN_0</ID>670 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add8</lparam></gate>
<gate>
<ID>360</ID>
<type>DA_FROM</type>
<position>68,-93</position>
<input>
<ID>IN_0</ID>451 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>215</ID>
<type>DA_FROM</type>
<position>-117.5,-135</position>
<input>
<ID>IN_0</ID>305 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo9</lparam></gate>
<gate>
<ID>546</ID>
<type>DA_FROM</type>
<position>-42,-192.5</position>
<input>
<ID>IN_0</ID>680 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>216</ID>
<type>DA_FROM</type>
<position>-108,-136</position>
<input>
<ID>IN_0</ID>297 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo10</lparam></gate>
<gate>
<ID>222</ID>
<type>DA_FROM</type>
<position>-117.5,-152</position>
<input>
<ID>IN_0</ID>304 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo13</lparam></gate>
<gate>
<ID>554</ID>
<type>FF_GND</type>
<position>27.5,-179.5</position>
<output>
<ID>OUT_0</ID>710 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>224</ID>
<type>DA_FROM</type>
<position>-108,-153</position>
<input>
<ID>IN_0</ID>295 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo14</lparam></gate>
<gate>
<ID>226</ID>
<type>DA_FROM</type>
<position>-117.5,-154</position>
<input>
<ID>IN_0</ID>303 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>258</ID>
<type>DE_TO</type>
<position>-16.5,-104</position>
<input>
<ID>IN_0</ID>331 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi0</lparam></gate>
<gate>
<ID>233</ID>
<type>DE_OR8</type>
<position>-23.5,-104</position>
<input>
<ID>IN_0</ID>414 </input>
<input>
<ID>IN_1</ID>325 </input>
<input>
<ID>IN_2</ID>334 </input>
<input>
<ID>IN_3</ID>335 </input>
<input>
<ID>IN_4</ID>346 </input>
<input>
<ID>IN_5</ID>343 </input>
<input>
<ID>IN_6</ID>341 </input>
<input>
<ID>IN_7</ID>338 </input>
<output>
<ID>OUT</ID>331 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>570</ID>
<type>AA_AND2</type>
<position>19,-188.5</position>
<input>
<ID>IN_0</ID>704 </input>
<input>
<ID>IN_1</ID>711 </input>
<output>
<ID>OUT</ID>703 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>-36,-89</position>
<input>
<ID>IN_0</ID>328 </input>
<input>
<ID>IN_1</ID>327 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AA_AND2</type>
<position>-50,-90</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>327 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>DA_FROM</type>
<position>-42,-88</position>
<input>
<ID>IN_0</ID>328 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>254</ID>
<type>DA_FROM</type>
<position>-58,-89</position>
<input>
<ID>IN_0</ID>329 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR0</lparam></gate>
<gate>
<ID>561</ID>
<type>DA_FROM</type>
<position>-3,-170.5</position>
<input>
<ID>IN_0</ID>693 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo9</lparam></gate>
<gate>
<ID>256</ID>
<type>DA_FROM</type>
<position>-58,-91</position>
<input>
<ID>IN_0</ID>330 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>565</ID>
<type>AA_AND2</type>
<position>19,-178.5</position>
<input>
<ID>IN_0</ID>699 </input>
<input>
<ID>IN_1</ID>692 </input>
<output>
<ID>OUT</ID>698 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>AA_AND2</type>
<position>-36,-94</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>333 </input>
<output>
<ID>OUT</ID>334 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>DA_FROM</type>
<position>-42,-93</position>
<input>
<ID>IN_0</ID>332 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>569</ID>
<type>DA_FROM</type>
<position>13,-182.5</position>
<input>
<ID>IN_0</ID>702 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>264</ID>
<type>DA_FROM</type>
<position>-42,-95</position>
<input>
<ID>IN_0</ID>333 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add0</lparam></gate>
<gate>
<ID>266</ID>
<type>AA_AND2</type>
<position>-36,-99</position>
<input>
<ID>IN_0</ID>336 </input>
<input>
<ID>IN_1</ID>329 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>573</ID>
<type>DA_FROM</type>
<position>13,-192.5</position>
<input>
<ID>IN_0</ID>706 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>268</ID>
<type>DA_FROM</type>
<position>-42,-98</position>
<input>
<ID>IN_0</ID>336 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>272</ID>
<type>AA_AND2</type>
<position>-36,-104</position>
<input>
<ID>IN_0</ID>340 </input>
<input>
<ID>IN_1</ID>339 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AE_SMALL_INVERTER</type>
<position>-51,-105</position>
<input>
<ID>IN_0</ID>330 </input>
<output>
<ID>OUT_0</ID>339 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>276</ID>
<type>DA_FROM</type>
<position>-42,-103</position>
<input>
<ID>IN_0</ID>340 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>-36,-109</position>
<input>
<ID>IN_0</ID>342 </input>
<input>
<ID>IN_1</ID>415 </input>
<output>
<ID>OUT</ID>341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>DA_FROM</type>
<position>-42,-108</position>
<input>
<ID>IN_0</ID>342 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>282</ID>
<type>AA_AND2</type>
<position>-36,-114</position>
<input>
<ID>IN_0</ID>344 </input>
<input>
<ID>IN_1</ID>416 </input>
<output>
<ID>OUT</ID>343 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>284</ID>
<type>DA_FROM</type>
<position>-42,-113</position>
<input>
<ID>IN_0</ID>344 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>286</ID>
<type>DA_FROM</type>
<position>-42,-118</position>
<input>
<ID>IN_0</ID>345 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_AND2</type>
<position>-36,-119</position>
<input>
<ID>IN_0</ID>345 </input>
<input>
<ID>IN_1</ID>347 </input>
<output>
<ID>OUT</ID>346 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>290</ID>
<type>DA_FROM</type>
<position>-42,-120</position>
<input>
<ID>IN_0</ID>347 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR0</lparam></gate>
<gate>
<ID>292</ID>
<type>DE_TO</type>
<position>-95,-158.5</position>
<input>
<ID>IN_0</ID>348 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>318</ID>
<type>DA_FROM</type>
<position>-42,-110</position>
<input>
<ID>IN_0</ID>415 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo1</lparam></gate>
<gate>
<ID>625</ID>
<type>DE_TO</type>
<position>148.5,-223</position>
<input>
<ID>IN_0</ID>772 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi15</lparam></gate>
<gate>
<ID>320</ID>
<type>DA_FROM</type>
<position>-42,-115</position>
<input>
<ID>IN_0</ID>416 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>629</ID>
<type>DA_FROM</type>
<position>123,-207</position>
<input>
<ID>IN_0</ID>769 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>324</ID>
<type>FF_GND</type>
<position>27.5,-100</position>
<output>
<ID>OUT_0</ID>440 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>660</ID>
<type>DA_FROM</type>
<position>68,-212</position>
<input>
<ID>IN_0</ID>799 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>325</ID>
<type>DE_TO</type>
<position>38.5,-104</position>
<input>
<ID>IN_0</ID>424 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi1</lparam></gate>
<gate>
<ID>326</ID>
<type>DE_OR8</type>
<position>31.5,-104</position>
<input>
<ID>IN_0</ID>440 </input>
<input>
<ID>IN_1</ID>419 </input>
<input>
<ID>IN_2</ID>427 </input>
<input>
<ID>IN_3</ID>428 </input>
<input>
<ID>IN_4</ID>438 </input>
<input>
<ID>IN_5</ID>435 </input>
<input>
<ID>IN_6</ID>433 </input>
<input>
<ID>IN_7</ID>430 </input>
<output>
<ID>OUT</ID>424 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>327</ID>
<type>AA_AND2</type>
<position>19,-89</position>
<input>
<ID>IN_0</ID>421 </input>
<input>
<ID>IN_1</ID>420 </input>
<output>
<ID>OUT</ID>419 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>633</ID>
<type>DA_FROM</type>
<position>123,-212</position>
<input>
<ID>IN_0</ID>773 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>5,-90</position>
<input>
<ID>IN_0</ID>422 </input>
<input>
<ID>IN_1</ID>423 </input>
<output>
<ID>OUT</ID>420 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>664</ID>
<type>AA_AND2</type>
<position>74,-223</position>
<input>
<ID>IN_0</ID>806 </input>
<input>
<ID>IN_1</ID>805 </input>
<output>
<ID>OUT</ID>804 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>DA_FROM</type>
<position>13,-88</position>
<input>
<ID>IN_0</ID>421 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>330</ID>
<type>DA_FROM</type>
<position>-3,-89</position>
<input>
<ID>IN_0</ID>422 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR1</lparam></gate>
<gate>
<ID>331</ID>
<type>DA_FROM</type>
<position>-3,-91</position>
<input>
<ID>IN_0</ID>423 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo1</lparam></gate>
<gate>
<ID>637</ID>
<type>AA_AND2</type>
<position>129,-223</position>
<input>
<ID>IN_0</ID>780 </input>
<input>
<ID>IN_1</ID>779 </input>
<output>
<ID>OUT</ID>778 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AA_AND2</type>
<position>19,-94</position>
<input>
<ID>IN_0</ID>425 </input>
<input>
<ID>IN_1</ID>426 </input>
<output>
<ID>OUT</ID>427 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>668</ID>
<type>AA_AND2</type>
<position>74,-233</position>
<input>
<ID>IN_0</ID>810 </input>
<input>
<ID>IN_1</ID>816 </input>
<output>
<ID>OUT</ID>809 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>DA_FROM</type>
<position>13,-93</position>
<input>
<ID>IN_0</ID>425 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>334</ID>
<type>DA_FROM</type>
<position>13,-95</position>
<input>
<ID>IN_0</ID>426 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add1</lparam></gate>
<gate>
<ID>335</ID>
<type>AA_AND2</type>
<position>19,-99</position>
<input>
<ID>IN_0</ID>429 </input>
<input>
<ID>IN_1</ID>422 </input>
<output>
<ID>OUT</ID>428 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>336</ID>
<type>DA_FROM</type>
<position>13,-98</position>
<input>
<ID>IN_0</ID>429 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>337</ID>
<type>AA_AND2</type>
<position>19,-104</position>
<input>
<ID>IN_0</ID>432 </input>
<input>
<ID>IN_1</ID>431 </input>
<output>
<ID>OUT</ID>430 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AE_SMALL_INVERTER</type>
<position>4,-105</position>
<input>
<ID>IN_0</ID>423 </input>
<output>
<ID>OUT_0</ID>431 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>339</ID>
<type>DA_FROM</type>
<position>13,-103</position>
<input>
<ID>IN_0</ID>432 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>517</ID>
<type>DA_FROM</type>
<position>68,-227</position>
<input>
<ID>IN_0</ID>808 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>19,-109</position>
<input>
<ID>IN_0</ID>434 </input>
<input>
<ID>IN_1</ID>441 </input>
<output>
<ID>OUT</ID>433 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>DA_FROM</type>
<position>13,-108</position>
<input>
<ID>IN_0</ID>434 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>342</ID>
<type>AA_AND2</type>
<position>19,-114</position>
<input>
<ID>IN_0</ID>436 </input>
<input>
<ID>IN_1</ID>442 </input>
<output>
<ID>OUT</ID>435 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>343</ID>
<type>DA_FROM</type>
<position>13,-113</position>
<input>
<ID>IN_0</ID>436 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>680</ID>
<type>AA_AND2</type>
<position>19,-208</position>
<input>
<ID>IN_0</ID>821 </input>
<input>
<ID>IN_1</ID>820 </input>
<output>
<ID>OUT</ID>819 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_AND2</type>
<position>19,-119</position>
<input>
<ID>IN_0</ID>437 </input>
<input>
<ID>IN_1</ID>439 </input>
<output>
<ID>OUT</ID>438 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>710</ID>
<type>AA_AND2</type>
<position>-36,-213</position>
<input>
<ID>IN_0</ID>851 </input>
<input>
<ID>IN_1</ID>852 </input>
<output>
<ID>OUT</ID>853 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>DA_FROM</type>
<position>13,-110</position>
<input>
<ID>IN_0</ID>441 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo2</lparam></gate>
<gate>
<ID>348</ID>
<type>DA_FROM</type>
<position>13,-115</position>
<input>
<ID>IN_0</ID>442 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>684</ID>
<type>AA_AND2</type>
<position>19,-213</position>
<input>
<ID>IN_0</ID>825 </input>
<input>
<ID>IN_1</ID>826 </input>
<output>
<ID>OUT</ID>827 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>351</ID>
<type>FF_GND</type>
<position>82.5,-100</position>
<output>
<ID>OUT_0</ID>466 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>688</ID>
<type>DA_FROM</type>
<position>13,-217</position>
<input>
<ID>IN_0</ID>829 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>353</ID>
<type>DE_OR8</type>
<position>86.5,-104</position>
<input>
<ID>IN_0</ID>466 </input>
<input>
<ID>IN_1</ID>445 </input>
<input>
<ID>IN_2</ID>453 </input>
<input>
<ID>IN_3</ID>454 </input>
<input>
<ID>IN_4</ID>464 </input>
<input>
<ID>IN_5</ID>461 </input>
<input>
<ID>IN_6</ID>459 </input>
<input>
<ID>IN_7</ID>456 </input>
<output>
<ID>OUT</ID>450 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>718</ID>
<type>AA_AND2</type>
<position>-36,-228</position>
<input>
<ID>IN_0</ID>860 </input>
<input>
<ID>IN_1</ID>867 </input>
<output>
<ID>OUT</ID>859 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>60,-90</position>
<input>
<ID>IN_0</ID>448 </input>
<input>
<ID>IN_1</ID>449 </input>
<output>
<ID>OUT</ID>446 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>692</ID>
<type>AA_AND2</type>
<position>19,-228</position>
<input>
<ID>IN_0</ID>834 </input>
<input>
<ID>IN_1</ID>841 </input>
<output>
<ID>OUT</ID>833 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>DA_FROM</type>
<position>52,-89</position>
<input>
<ID>IN_0</ID>448 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR2</lparam></gate>
<gate>
<ID>358</ID>
<type>DA_FROM</type>
<position>52,-91</position>
<input>
<ID>IN_0</ID>449 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo2</lparam></gate>
<gate>
<ID>706</ID>
<type>AA_AND2</type>
<position>-50,-209</position>
<input>
<ID>IN_0</ID>848 </input>
<input>
<ID>IN_1</ID>849 </input>
<output>
<ID>OUT</ID>846 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>74,-94</position>
<input>
<ID>IN_0</ID>451 </input>
<input>
<ID>IN_1</ID>452 </input>
<output>
<ID>OUT</ID>453 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>361</ID>
<type>DA_FROM</type>
<position>68,-95</position>
<input>
<ID>IN_0</ID>452 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add2</lparam></gate>
<gate>
<ID>726</ID>
<type>DA_FROM</type>
<position>-42,-234</position>
<input>
<ID>IN_0</ID>868 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo11</lparam></gate>
<gate>
<ID>363</ID>
<type>DA_FROM</type>
<position>68,-98</position>
<input>
<ID>IN_0</ID>455 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>700</ID>
<type>DA_FROM</type>
<position>13,-234</position>
<input>
<ID>IN_0</ID>842 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo12</lparam></gate>
<gate>
<ID>365</ID>
<type>AE_SMALL_INVERTER</type>
<position>59,-105</position>
<input>
<ID>IN_0</ID>449 </input>
<output>
<ID>OUT_0</ID>457 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>714</ID>
<type>DA_FROM</type>
<position>-42,-217</position>
<input>
<ID>IN_0</ID>855 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>367</ID>
<type>AA_AND2</type>
<position>74,-109</position>
<input>
<ID>IN_0</ID>460 </input>
<input>
<ID>IN_1</ID>467 </input>
<output>
<ID>OUT</ID>459 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>545</ID>
<type>AA_AND2</type>
<position>-36,-193.5</position>
<input>
<ID>IN_0</ID>680 </input>
<input>
<ID>IN_1</ID>686 </input>
<output>
<ID>OUT</ID>679 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>368</ID>
<type>DA_FROM</type>
<position>68,-108</position>
<input>
<ID>IN_0</ID>460 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>576</ID>
<type>DA_FROM</type>
<position>13,-194.5</position>
<input>
<ID>IN_0</ID>712 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo8</lparam></gate>
<gate>
<ID>369</ID>
<type>AA_AND2</type>
<position>74,-114</position>
<input>
<ID>IN_0</ID>462 </input>
<input>
<ID>IN_1</ID>468 </input>
<output>
<ID>OUT</ID>461 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>370</ID>
<type>DA_FROM</type>
<position>68,-113</position>
<input>
<ID>IN_0</ID>462 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>734</ID>
<type>FF_GND</type>
<position>82.5,-189</position>
<output>
<ID>OUT_0</ID>873 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>371</ID>
<type>DA_FROM</type>
<position>68,-118</position>
<input>
<ID>IN_0</ID>463 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>580</ID>
<type>AA_AND2</type>
<position>60,-169.5</position>
<input>
<ID>IN_0</ID>718 </input>
<input>
<ID>IN_1</ID>719 </input>
<output>
<ID>OUT</ID>716 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>373</ID>
<type>DA_FROM</type>
<position>68,-120</position>
<input>
<ID>IN_0</ID>465 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR2</lparam></gate>
<gate>
<ID>374</ID>
<type>DA_FROM</type>
<position>68,-110</position>
<input>
<ID>IN_0</ID>467 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo3</lparam></gate>
<gate>
<ID>375</ID>
<type>DA_FROM</type>
<position>68,-115</position>
<input>
<ID>IN_0</ID>468 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo1</lparam></gate>
<gate>
<ID>584</ID>
<type>DA_FROM</type>
<position>68,-174.5</position>
<input>
<ID>IN_0</ID>722 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add10</lparam></gate>
<gate>
<ID>378</ID>
<type>FF_GND</type>
<position>137.5,-100</position>
<output>
<ID>OUT_0</ID>496 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>742</ID>
<type>FF_GND</type>
<position>82.5,-228.5</position>
<output>
<ID>OUT_0</ID>877 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>379</ID>
<type>DE_TO</type>
<position>148.5,-104</position>
<input>
<ID>IN_0</ID>476 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi3</lparam></gate>
<gate>
<ID>557</ID>
<type>AA_AND2</type>
<position>19,-168.5</position>
<input>
<ID>IN_0</ID>691 </input>
<input>
<ID>IN_1</ID>690 </input>
<output>
<ID>OUT</ID>689 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>380</ID>
<type>DE_OR8</type>
<position>141.5,-104</position>
<input>
<ID>IN_0</ID>496 </input>
<input>
<ID>IN_1</ID>471 </input>
<input>
<ID>IN_2</ID>479 </input>
<input>
<ID>IN_3</ID>480 </input>
<input>
<ID>IN_4</ID>494 </input>
<input>
<ID>IN_5</ID>491 </input>
<input>
<ID>IN_6</ID>485 </input>
<input>
<ID>IN_7</ID>482 </input>
<output>
<ID>OUT</ID>476 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>588</ID>
<type>DA_FROM</type>
<position>68,-187.5</position>
<input>
<ID>IN_0</ID>730 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>381</ID>
<type>AA_AND2</type>
<position>129,-89</position>
<input>
<ID>IN_0</ID>473 </input>
<input>
<ID>IN_1</ID>472 </input>
<output>
<ID>OUT</ID>471 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>382</ID>
<type>AA_AND2</type>
<position>115,-90</position>
<input>
<ID>IN_0</ID>474 </input>
<input>
<ID>IN_1</ID>475 </input>
<output>
<ID>OUT</ID>472 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>730</ID>
<type>FF_GND</type>
<position>-27.5,-189</position>
<output>
<ID>OUT_0</ID>871 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>383</ID>
<type>DA_FROM</type>
<position>123,-88</position>
<input>
<ID>IN_0</ID>473 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>689</ID>
<type>AA_AND2</type>
<position>19,-223</position>
<input>
<ID>IN_0</ID>832 </input>
<input>
<ID>IN_1</ID>831 </input>
<output>
<ID>OUT</ID>830 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>384</ID>
<type>DA_FROM</type>
<position>107,-89</position>
<input>
<ID>IN_0</ID>474 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR3</lparam></gate>
<gate>
<ID>720</ID>
<type>AA_AND2</type>
<position>-36,-233</position>
<input>
<ID>IN_0</ID>862 </input>
<input>
<ID>IN_1</ID>868 </input>
<output>
<ID>OUT</ID>861 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>385</ID>
<type>DA_FROM</type>
<position>107,-91</position>
<input>
<ID>IN_0</ID>475 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo3</lparam></gate>
<gate>
<ID>551</ID>
<type>DA_FROM</type>
<position>-42,-194.5</position>
<input>
<ID>IN_0</ID>686 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo7</lparam></gate>
<gate>
<ID>386</ID>
<type>AA_AND2</type>
<position>129,-94</position>
<input>
<ID>IN_0</ID>477 </input>
<input>
<ID>IN_1</ID>478 </input>
<output>
<ID>OUT</ID>479 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>387</ID>
<type>DA_FROM</type>
<position>123,-93</position>
<input>
<ID>IN_0</ID>477 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>693</ID>
<type>DA_FROM</type>
<position>13,-227</position>
<input>
<ID>IN_0</ID>834 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>388</ID>
<type>DA_FROM</type>
<position>123,-95</position>
<input>
<ID>IN_0</ID>478 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add3</lparam></gate>
<gate>
<ID>389</ID>
<type>AA_AND2</type>
<position>129,-99</position>
<input>
<ID>IN_0</ID>481 </input>
<input>
<ID>IN_1</ID>474 </input>
<output>
<ID>OUT</ID>480 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>539</ID>
<type>DA_FROM</type>
<position>-42,-177.5</position>
<input>
<ID>IN_0</ID>673 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>390</ID>
<type>DA_FROM</type>
<position>123,-98</position>
<input>
<ID>IN_0</ID>481 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>391</ID>
<type>AA_AND2</type>
<position>129,-104</position>
<input>
<ID>IN_0</ID>484 </input>
<input>
<ID>IN_1</ID>483 </input>
<output>
<ID>OUT</ID>482 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>392</ID>
<type>AE_SMALL_INVERTER</type>
<position>114,-105</position>
<input>
<ID>IN_0</ID>475 </input>
<output>
<ID>OUT_0</ID>483 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>393</ID>
<type>DA_FROM</type>
<position>123,-103</position>
<input>
<ID>IN_0</ID>484 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>559</ID>
<type>DA_FROM</type>
<position>13,-167.5</position>
<input>
<ID>IN_0</ID>691 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>394</ID>
<type>AA_AND2</type>
<position>129,-109</position>
<input>
<ID>IN_0</ID>490 </input>
<input>
<ID>IN_1</ID>497 </input>
<output>
<ID>OUT</ID>485 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>395</ID>
<type>DA_FROM</type>
<position>123,-108</position>
<input>
<ID>IN_0</ID>490 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>396</ID>
<type>AA_AND2</type>
<position>129,-114</position>
<input>
<ID>IN_0</ID>492 </input>
<input>
<ID>IN_1</ID>498 </input>
<output>
<ID>OUT</ID>491 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>732</ID>
<type>FF_GND</type>
<position>27.5,-189</position>
<output>
<ID>OUT_0</ID>872 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>397</ID>
<type>DA_FROM</type>
<position>123,-113</position>
<input>
<ID>IN_0</ID>492 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>398</ID>
<type>DA_FROM</type>
<position>123,-118</position>
<input>
<ID>IN_0</ID>493 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>399</ID>
<type>AA_AND2</type>
<position>129,-119</position>
<input>
<ID>IN_0</ID>493 </input>
<input>
<ID>IN_1</ID>495 </input>
<output>
<ID>OUT</ID>494 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>400</ID>
<type>DA_FROM</type>
<position>123,-120</position>
<input>
<ID>IN_0</ID>495 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR3</lparam></gate>
<gate>
<ID>736</ID>
<type>FF_GND</type>
<position>137.5,-189</position>
<output>
<ID>OUT_0</ID>874 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>401</ID>
<type>DA_FROM</type>
<position>123,-110</position>
<input>
<ID>IN_0</ID>497 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo4</lparam></gate>
<gate>
<ID>567</ID>
<type>AA_AND2</type>
<position>19,-183.5</position>
<input>
<ID>IN_0</ID>702 </input>
<input>
<ID>IN_1</ID>701 </input>
<output>
<ID>OUT</ID>700 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>402</ID>
<type>DA_FROM</type>
<position>123,-115</position>
<input>
<ID>IN_0</ID>498 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo2</lparam></gate>
<gate>
<ID>581</ID>
<type>DA_FROM</type>
<position>52,-168.5</position>
<input>
<ID>IN_0</ID>718 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR10</lparam></gate>
<gate>
<ID>740</ID>
<type>FF_GND</type>
<position>27.5,-228.5</position>
<output>
<ID>OUT_0</ID>876 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>405</ID>
<type>FF_GND</type>
<position>137.5,-139.5</position>
<output>
<ID>OUT_0</ID>531 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>555</ID>
<type>DE_TO</type>
<position>38.5,-183.5</position>
<input>
<ID>IN_0</ID>694 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi9</lparam></gate>
<gate>
<ID>406</ID>
<type>DE_TO</type>
<position>148.5,-143.5</position>
<input>
<ID>IN_0</ID>506 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi7</lparam></gate>
<gate>
<ID>407</ID>
<type>DE_OR8</type>
<position>141.5,-143.5</position>
<input>
<ID>IN_0</ID>531 </input>
<input>
<ID>IN_1</ID>501 </input>
<input>
<ID>IN_2</ID>509 </input>
<input>
<ID>IN_3</ID>510 </input>
<input>
<ID>IN_4</ID>529 </input>
<input>
<ID>IN_5</ID>526 </input>
<input>
<ID>IN_6</ID>524 </input>
<input>
<ID>IN_7</ID>512 </input>
<output>
<ID>OUT</ID>506 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>585</ID>
<type>DA_FROM</type>
<position>68,-177.5</position>
<input>
<ID>IN_0</ID>725 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>408</ID>
<type>AA_AND2</type>
<position>129,-128.5</position>
<input>
<ID>IN_0</ID>503 </input>
<input>
<ID>IN_1</ID>502 </input>
<output>
<ID>OUT</ID>501 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>744</ID>
<type>FF_GND</type>
<position>137.5,-228.5</position>
<output>
<ID>OUT_0</ID>878 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>409</ID>
<type>AA_AND2</type>
<position>115,-129.5</position>
<input>
<ID>IN_0</ID>504 </input>
<input>
<ID>IN_1</ID>505 </input>
<output>
<ID>OUT</ID>502 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>575</ID>
<type>DA_FROM</type>
<position>13,-189.5</position>
<input>
<ID>IN_0</ID>711 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo10</lparam></gate>
<gate>
<ID>410</ID>
<type>DA_FROM</type>
<position>123,-127.5</position>
<input>
<ID>IN_0</ID>503 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>411</ID>
<type>DA_FROM</type>
<position>107,-128.5</position>
<input>
<ID>IN_0</ID>504 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR7</lparam></gate>
<gate>
<ID>589</ID>
<type>AA_AND2</type>
<position>74,-193.5</position>
<input>
<ID>IN_0</ID>732 </input>
<input>
<ID>IN_1</ID>738 </input>
<output>
<ID>OUT</ID>731 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>412</ID>
<type>DA_FROM</type>
<position>107,-130.5</position>
<input>
<ID>IN_0</ID>505 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo7</lparam></gate>
<gate>
<ID>413</ID>
<type>AA_AND2</type>
<position>129,-133.5</position>
<input>
<ID>IN_0</ID>507 </input>
<input>
<ID>IN_1</ID>508 </input>
<output>
<ID>OUT</ID>509 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>563</ID>
<type>DA_FROM</type>
<position>13,-172.5</position>
<input>
<ID>IN_0</ID>695 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>414</ID>
<type>DA_FROM</type>
<position>123,-132.5</position>
<input>
<ID>IN_0</ID>507 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>415</ID>
<type>DA_FROM</type>
<position>123,-134.5</position>
<input>
<ID>IN_0</ID>508 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add7</lparam></gate>
<gate>
<ID>593</ID>
<type>DA_FROM</type>
<position>68,-189.5</position>
<input>
<ID>IN_0</ID>737 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo11</lparam></gate>
<gate>
<ID>416</ID>
<type>AA_AND2</type>
<position>129,-138.5</position>
<input>
<ID>IN_0</ID>511 </input>
<input>
<ID>IN_1</ID>504 </input>
<output>
<ID>OUT</ID>510 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>417</ID>
<type>DA_FROM</type>
<position>123,-137.5</position>
<input>
<ID>IN_0</ID>511 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>418</ID>
<type>AA_AND2</type>
<position>129,-143.5</position>
<input>
<ID>IN_0</ID>523 </input>
<input>
<ID>IN_1</ID>522 </input>
<output>
<ID>OUT</ID>512 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>419</ID>
<type>AE_SMALL_INVERTER</type>
<position>114,-144.5</position>
<input>
<ID>IN_0</ID>505 </input>
<output>
<ID>OUT_0</ID>522 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>597</ID>
<type>FF_GND</type>
<position>137.5,-179.5</position>
<output>
<ID>OUT_0</ID>762 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>420</ID>
<type>DA_FROM</type>
<position>123,-142.5</position>
<input>
<ID>IN_0</ID>523 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>421</ID>
<type>AA_AND2</type>
<position>129,-148.5</position>
<input>
<ID>IN_0</ID>525 </input>
<input>
<ID>IN_1</ID>532 </input>
<output>
<ID>OUT</ID>524 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>571</ID>
<type>DA_FROM</type>
<position>13,-187.5</position>
<input>
<ID>IN_0</ID>704 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>422</ID>
<type>DA_FROM</type>
<position>123,-147.5</position>
<input>
<ID>IN_0</ID>525 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>423</ID>
<type>AA_AND2</type>
<position>129,-153.5</position>
<input>
<ID>IN_0</ID>527 </input>
<input>
<ID>IN_1</ID>533 </input>
<output>
<ID>OUT</ID>526 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>601</ID>
<type>AA_AND2</type>
<position>115,-169.5</position>
<input>
<ID>IN_0</ID>744 </input>
<input>
<ID>IN_1</ID>745 </input>
<output>
<ID>OUT</ID>742 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>424</ID>
<type>DA_FROM</type>
<position>123,-152.5</position>
<input>
<ID>IN_0</ID>527 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>425</ID>
<type>DA_FROM</type>
<position>123,-157.5</position>
<input>
<ID>IN_0</ID>528 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>426</ID>
<type>AA_AND2</type>
<position>129,-158.5</position>
<input>
<ID>IN_0</ID>528 </input>
<input>
<ID>IN_1</ID>530 </input>
<output>
<ID>OUT</ID>529 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>427</ID>
<type>DA_FROM</type>
<position>123,-159.5</position>
<input>
<ID>IN_0</ID>530 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR7</lparam></gate>
<gate>
<ID>605</ID>
<type>AA_AND2</type>
<position>129,-173.5</position>
<input>
<ID>IN_0</ID>747 </input>
<input>
<ID>IN_1</ID>748 </input>
<output>
<ID>OUT</ID>749 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>428</ID>
<type>DA_FROM</type>
<position>123,-149.5</position>
<input>
<ID>IN_0</ID>532 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo8</lparam></gate>
<gate>
<ID>429</ID>
<type>DA_FROM</type>
<position>123,-154.5</position>
<input>
<ID>IN_0</ID>533 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo6</lparam></gate>
<gate>
<ID>609</ID>
<type>DA_FROM</type>
<position>123,-177.5</position>
<input>
<ID>IN_0</ID>751 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>432</ID>
<type>FF_GND</type>
<position>82.5,-139.5</position>
<output>
<ID>OUT_0</ID>606 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>640</ID>
<type>AA_AND2</type>
<position>129,-228</position>
<input>
<ID>IN_0</ID>782 </input>
<input>
<ID>IN_1</ID>789 </input>
<output>
<ID>OUT</ID>781 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>433</ID>
<type>DE_TO</type>
<position>93.5,-143.5</position>
<input>
<ID>IN_0</ID>541 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi6</lparam></gate>
<gate>
<ID>434</ID>
<type>DE_OR8</type>
<position>86.5,-143.5</position>
<input>
<ID>IN_0</ID>606 </input>
<input>
<ID>IN_1</ID>536 </input>
<input>
<ID>IN_2</ID>586 </input>
<input>
<ID>IN_3</ID>587 </input>
<input>
<ID>IN_4</ID>604 </input>
<input>
<ID>IN_5</ID>601 </input>
<input>
<ID>IN_6</ID>599 </input>
<input>
<ID>IN_7</ID>589 </input>
<output>
<ID>OUT</ID>541 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>435</ID>
<type>AA_AND2</type>
<position>74,-128.5</position>
<input>
<ID>IN_0</ID>538 </input>
<input>
<ID>IN_1</ID>537 </input>
<output>
<ID>OUT</ID>536 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>613</ID>
<type>AA_AND2</type>
<position>129,-188.5</position>
<input>
<ID>IN_0</ID>756 </input>
<input>
<ID>IN_1</ID>763 </input>
<output>
<ID>OUT</ID>755 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>436</ID>
<type>AA_AND2</type>
<position>60,-129.5</position>
<input>
<ID>IN_0</ID>539 </input>
<input>
<ID>IN_1</ID>540 </input>
<output>
<ID>OUT</ID>537 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>437</ID>
<type>DA_FROM</type>
<position>68,-127.5</position>
<input>
<ID>IN_0</ID>538 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>438</ID>
<type>DA_FROM</type>
<position>52,-128.5</position>
<input>
<ID>IN_0</ID>539 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR6</lparam></gate>
<gate>
<ID>439</ID>
<type>DA_FROM</type>
<position>52,-130.5</position>
<input>
<ID>IN_0</ID>540 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo6</lparam></gate>
<gate>
<ID>440</ID>
<type>AA_AND2</type>
<position>74,-133.5</position>
<input>
<ID>IN_0</ID>579 </input>
<input>
<ID>IN_1</ID>585 </input>
<output>
<ID>OUT</ID>586 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>648</ID>
<type>DA_FROM</type>
<position>123,-234</position>
<input>
<ID>IN_0</ID>790 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo14</lparam></gate>
<gate>
<ID>441</ID>
<type>DA_FROM</type>
<position>68,-132.5</position>
<input>
<ID>IN_0</ID>579 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>442</ID>
<type>DA_FROM</type>
<position>68,-134.5</position>
<input>
<ID>IN_0</ID>585 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add6</lparam></gate>
<gate>
<ID>443</ID>
<type>AA_AND2</type>
<position>74,-138.5</position>
<input>
<ID>IN_0</ID>588 </input>
<input>
<ID>IN_1</ID>539 </input>
<output>
<ID>OUT</ID>587 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>621</ID>
<type>DA_FROM</type>
<position>123,-194.5</position>
<input>
<ID>IN_0</ID>764 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo10</lparam></gate>
<gate>
<ID>444</ID>
<type>DA_FROM</type>
<position>68,-137.5</position>
<input>
<ID>IN_0</ID>588 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>652</ID>
<type>DE_TO</type>
<position>93.5,-223</position>
<input>
<ID>IN_0</ID>798 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi14</lparam></gate>
<gate>
<ID>445</ID>
<type>AA_AND2</type>
<position>74,-143.5</position>
<input>
<ID>IN_0</ID>598 </input>
<input>
<ID>IN_1</ID>590 </input>
<output>
<ID>OUT</ID>589 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>446</ID>
<type>AE_SMALL_INVERTER</type>
<position>59,-144.5</position>
<input>
<ID>IN_0</ID>540 </input>
<output>
<ID>OUT_0</ID>590 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>447</ID>
<type>DA_FROM</type>
<position>68,-142.5</position>
<input>
<ID>IN_0</ID>598 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>448</ID>
<type>AA_AND2</type>
<position>74,-148.5</position>
<input>
<ID>IN_0</ID>600 </input>
<input>
<ID>IN_1</ID>607 </input>
<output>
<ID>OUT</ID>599 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>615</ID>
<type>AA_AND2</type>
<position>129,-193.5</position>
<input>
<ID>IN_0</ID>758 </input>
<input>
<ID>IN_1</ID>764 </input>
<output>
<ID>OUT</ID>757 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>450</ID>
<type>AA_AND2</type>
<position>74,-153.5</position>
<input>
<ID>IN_0</ID>602 </input>
<input>
<ID>IN_1</ID>608 </input>
<output>
<ID>OUT</ID>601 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>451</ID>
<type>DA_FROM</type>
<position>68,-152.5</position>
<input>
<ID>IN_0</ID>602 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>452</ID>
<type>DA_FROM</type>
<position>68,-157.5</position>
<input>
<ID>IN_0</ID>603 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>453</ID>
<type>AA_AND2</type>
<position>74,-158.5</position>
<input>
<ID>IN_0</ID>603 </input>
<input>
<ID>IN_1</ID>605 </input>
<output>
<ID>OUT</ID>604 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>603</ID>
<type>DA_FROM</type>
<position>107,-168.5</position>
<input>
<ID>IN_0</ID>744 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR11</lparam></gate>
<gate>
<ID>454</ID>
<type>DA_FROM</type>
<position>68,-159.5</position>
<input>
<ID>IN_0</ID>605 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR6</lparam></gate>
<gate>
<ID>455</ID>
<type>DA_FROM</type>
<position>68,-149.5</position>
<input>
<ID>IN_0</ID>607 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo7</lparam></gate>
<gate>
<ID>456</ID>
<type>DA_FROM</type>
<position>68,-154.5</position>
<input>
<ID>IN_0</ID>608 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo5</lparam></gate>
<gate>
<ID>459</ID>
<type>FF_GND</type>
<position>27.5,-139.5</position>
<output>
<ID>OUT_0</ID>632 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>460</ID>
<type>DE_TO</type>
<position>38.5,-143.5</position>
<input>
<ID>IN_0</ID>616 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi5</lparam></gate>
<gate>
<ID>461</ID>
<type>DE_OR8</type>
<position>31.5,-143.5</position>
<input>
<ID>IN_0</ID>632 </input>
<input>
<ID>IN_1</ID>611 </input>
<input>
<ID>IN_2</ID>619 </input>
<input>
<ID>IN_3</ID>620 </input>
<input>
<ID>IN_4</ID>630 </input>
<input>
<ID>IN_5</ID>627 </input>
<input>
<ID>IN_6</ID>625 </input>
<input>
<ID>IN_7</ID>622 </input>
<output>
<ID>OUT</ID>616 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>611</ID>
<type>AE_SMALL_INVERTER</type>
<position>114,-184.5</position>
<input>
<ID>IN_0</ID>745 </input>
<output>
<ID>OUT_0</ID>753 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>462</ID>
<type>AA_AND2</type>
<position>19,-128.5</position>
<input>
<ID>IN_0</ID>613 </input>
<input>
<ID>IN_1</ID>612 </input>
<output>
<ID>OUT</ID>611 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>463</ID>
<type>AA_AND2</type>
<position>5,-129.5</position>
<input>
<ID>IN_0</ID>614 </input>
<input>
<ID>IN_1</ID>615 </input>
<output>
<ID>OUT</ID>612 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>641</ID>
<type>DA_FROM</type>
<position>123,-227</position>
<input>
<ID>IN_0</ID>782 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>464</ID>
<type>DA_FROM</type>
<position>13,-127.5</position>
<input>
<ID>IN_0</ID>613 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>631</ID>
<type>DA_FROM</type>
<position>107,-210</position>
<input>
<ID>IN_0</ID>771 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>466</ID>
<type>DA_FROM</type>
<position>-3,-130.5</position>
<input>
<ID>IN_0</ID>615 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo5</lparam></gate>
<gate>
<ID>467</ID>
<type>AA_AND2</type>
<position>19,-133.5</position>
<input>
<ID>IN_0</ID>617 </input>
<input>
<ID>IN_1</ID>618 </input>
<output>
<ID>OUT</ID>619 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>468</ID>
<type>DA_FROM</type>
<position>13,-132.5</position>
<input>
<ID>IN_0</ID>617 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>469</ID>
<type>DA_FROM</type>
<position>13,-134.5</position>
<input>
<ID>IN_0</ID>618 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add5</lparam></gate>
<gate>
<ID>470</ID>
<type>AA_AND2</type>
<position>19,-138.5</position>
<input>
<ID>IN_0</ID>621 </input>
<input>
<ID>IN_1</ID>614 </input>
<output>
<ID>OUT</ID>620 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>471</ID>
<type>DA_FROM</type>
<position>13,-137.5</position>
<input>
<ID>IN_0</ID>621 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>472</ID>
<type>AA_AND2</type>
<position>19,-143.5</position>
<input>
<ID>IN_0</ID>624 </input>
<input>
<ID>IN_1</ID>623 </input>
<output>
<ID>OUT</ID>622 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>473</ID>
<type>AE_SMALL_INVERTER</type>
<position>4,-144.5</position>
<input>
<ID>IN_0</ID>615 </input>
<output>
<ID>OUT_0</ID>623 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>639</ID>
<type>DA_FROM</type>
<position>123,-222</position>
<input>
<ID>IN_0</ID>780 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>474</ID>
<type>DA_FROM</type>
<position>13,-142.5</position>
<input>
<ID>IN_0</ID>624 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>475</ID>
<type>AA_AND2</type>
<position>19,-148.5</position>
<input>
<ID>IN_0</ID>626 </input>
<input>
<ID>IN_1</ID>633 </input>
<output>
<ID>OUT</ID>625 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>653</ID>
<type>DE_OR8</type>
<position>86.5,-223</position>
<input>
<ID>IN_0</ID>814 </input>
<input>
<ID>IN_1</ID>793 </input>
<input>
<ID>IN_2</ID>801 </input>
<input>
<ID>IN_3</ID>802 </input>
<input>
<ID>IN_4</ID>877 </input>
<input>
<ID>IN_5</ID>809 </input>
<input>
<ID>IN_6</ID>807 </input>
<input>
<ID>IN_7</ID>804 </input>
<output>
<ID>OUT</ID>798 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>476</ID>
<type>DA_FROM</type>
<position>13,-147.5</position>
<input>
<ID>IN_0</ID>626 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>477</ID>
<type>AA_AND2</type>
<position>19,-153.5</position>
<input>
<ID>IN_0</ID>628 </input>
<input>
<ID>IN_1</ID>634 </input>
<output>
<ID>OUT</ID>627 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>627</ID>
<type>AA_AND2</type>
<position>129,-208</position>
<input>
<ID>IN_0</ID>769 </input>
<input>
<ID>IN_1</ID>768 </input>
<output>
<ID>OUT</ID>767 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>478</ID>
<type>DA_FROM</type>
<position>13,-152.5</position>
<input>
<ID>IN_0</ID>628 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>479</ID>
<type>DA_FROM</type>
<position>13,-157.5</position>
<input>
<ID>IN_0</ID>629 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>657</ID>
<type>DA_FROM</type>
<position>52,-208</position>
<input>
<ID>IN_0</ID>796 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR14</lparam></gate>
<gate>
<ID>480</ID>
<type>AA_AND2</type>
<position>19,-158.5</position>
<input>
<ID>IN_0</ID>629 </input>
<input>
<ID>IN_1</ID>631 </input>
<output>
<ID>OUT</ID>630 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>481</ID>
<type>DA_FROM</type>
<position>13,-159.5</position>
<input>
<ID>IN_0</ID>631 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR5</lparam></gate>
<gate>
<ID>482</ID>
<type>DA_FROM</type>
<position>13,-149.5</position>
<input>
<ID>IN_0</ID>633 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo6</lparam></gate>
<gate>
<ID>483</ID>
<type>DA_FROM</type>
<position>13,-154.5</position>
<input>
<ID>IN_0</ID>634 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo4</lparam></gate>
<gate>
<ID>661</ID>
<type>DA_FROM</type>
<position>68,-214</position>
<input>
<ID>IN_0</ID>800 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add14</lparam></gate>
<gate>
<ID>635</ID>
<type>AA_AND2</type>
<position>129,-218</position>
<input>
<ID>IN_0</ID>777 </input>
<input>
<ID>IN_1</ID>770 </input>
<output>
<ID>OUT</ID>776 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>486</ID>
<type>FF_GND</type>
<position>-27.5,-139.5</position>
<output>
<ID>OUT_0</ID>658 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>487</ID>
<type>DE_TO</type>
<position>-16.5,-143.5</position>
<input>
<ID>IN_0</ID>642 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi4</lparam></gate>
<gate>
<ID>665</ID>
<type>AE_SMALL_INVERTER</type>
<position>59,-224</position>
<input>
<ID>IN_0</ID>797 </input>
<output>
<ID>OUT_0</ID>805 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>488</ID>
<type>DE_OR8</type>
<position>-23.5,-143.5</position>
<input>
<ID>IN_0</ID>658 </input>
<input>
<ID>IN_1</ID>637 </input>
<input>
<ID>IN_2</ID>645 </input>
<input>
<ID>IN_3</ID>646 </input>
<input>
<ID>IN_4</ID>656 </input>
<input>
<ID>IN_5</ID>653 </input>
<input>
<ID>IN_6</ID>651 </input>
<input>
<ID>IN_7</ID>648 </input>
<output>
<ID>OUT</ID>642 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>489</ID>
<type>AA_AND2</type>
<position>-36,-128.5</position>
<input>
<ID>IN_0</ID>639 </input>
<input>
<ID>IN_1</ID>638 </input>
<output>
<ID>OUT</ID>637 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>527</ID>
<type>DA_FROM</type>
<position>68,-172.5</position>
<input>
<ID>IN_0</ID>721 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>490</ID>
<type>AA_AND2</type>
<position>-50,-129.5</position>
<input>
<ID>IN_0</ID>640 </input>
<input>
<ID>IN_1</ID>641 </input>
<output>
<ID>OUT</ID>638 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>491</ID>
<type>DA_FROM</type>
<position>-42,-127.5</position>
<input>
<ID>IN_0</ID>639 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>669</ID>
<type>DA_FROM</type>
<position>68,-232</position>
<input>
<ID>IN_0</ID>810 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>492</ID>
<type>DA_FROM</type>
<position>-58,-128.5</position>
<input>
<ID>IN_0</ID>640 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR4</lparam></gate>
<gate>
<ID>493</ID>
<type>DA_FROM</type>
<position>-58,-130.5</position>
<input>
<ID>IN_0</ID>641 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo4</lparam></gate>
<gate>
<ID>494</ID>
<type>AA_AND2</type>
<position>-36,-133.5</position>
<input>
<ID>IN_0</ID>643 </input>
<input>
<ID>IN_1</ID>644 </input>
<output>
<ID>OUT</ID>645 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>495</ID>
<type>DA_FROM</type>
<position>-42,-132.5</position>
<input>
<ID>IN_0</ID>643 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>673</ID>
<type>DA_FROM</type>
<position>68,-229</position>
<input>
<ID>IN_0</ID>815 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>496</ID>
<type>DA_FROM</type>
<position>-42,-134.5</position>
<input>
<ID>IN_0</ID>644 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add4</lparam></gate>
<gate>
<ID>704</ID>
<type>DE_OR8</type>
<position>-23.5,-223</position>
<input>
<ID>IN_0</ID>866 </input>
<input>
<ID>IN_1</ID>845 </input>
<input>
<ID>IN_2</ID>853 </input>
<input>
<ID>IN_3</ID>854 </input>
<input>
<ID>IN_4</ID>875 </input>
<input>
<ID>IN_5</ID>861 </input>
<input>
<ID>IN_6</ID>859 </input>
<input>
<ID>IN_7</ID>856 </input>
<output>
<ID>OUT</ID>850 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>497</ID>
<type>AA_AND2</type>
<position>-36,-138.5</position>
<input>
<ID>IN_0</ID>647 </input>
<input>
<ID>IN_1</ID>640 </input>
<output>
<ID>OUT</ID>646 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>535</ID>
<type>AA_AND2</type>
<position>-36,-173.5</position>
<input>
<ID>IN_0</ID>669 </input>
<input>
<ID>IN_1</ID>670 </input>
<output>
<ID>OUT</ID>671 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>498</ID>
<type>DA_FROM</type>
<position>-42,-137.5</position>
<input>
<ID>IN_0</ID>647 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>499</ID>
<type>AA_AND2</type>
<position>-36,-143.5</position>
<input>
<ID>IN_0</ID>650 </input>
<input>
<ID>IN_1</ID>649 </input>
<output>
<ID>OUT</ID>648 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>677</ID>
<type>FF_GND</type>
<position>27.5,-219</position>
<output>
<ID>OUT_0</ID>840 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>500</ID>
<type>AE_SMALL_INVERTER</type>
<position>-51,-144.5</position>
<input>
<ID>IN_0</ID>641 </input>
<output>
<ID>OUT_0</ID>649 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>708</ID>
<type>DA_FROM</type>
<position>-58,-208</position>
<input>
<ID>IN_0</ID>848 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR12</lparam></gate>
<gate>
<ID>501</ID>
<type>DA_FROM</type>
<position>-42,-142.5</position>
<input>
<ID>IN_0</ID>650 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>523</ID>
<type>DE_TO</type>
<position>93.5,-183.5</position>
<input>
<ID>IN_0</ID>720 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi10</lparam></gate>
<gate>
<ID>502</ID>
<type>AA_AND2</type>
<position>-36,-148.5</position>
<input>
<ID>IN_0</ID>652 </input>
<input>
<ID>IN_1</ID>659 </input>
<output>
<ID>OUT</ID>651 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>503</ID>
<type>DA_FROM</type>
<position>-42,-147.5</position>
<input>
<ID>IN_0</ID>652 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>681</ID>
<type>AA_AND2</type>
<position>5,-209</position>
<input>
<ID>IN_0</ID>822 </input>
<input>
<ID>IN_1</ID>823 </input>
<output>
<ID>OUT</ID>820 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>504</ID>
<type>AA_AND2</type>
<position>-36,-153.5</position>
<input>
<ID>IN_0</ID>654 </input>
<input>
<ID>IN_1</ID>660 </input>
<output>
<ID>OUT</ID>653 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>712</ID>
<type>DA_FROM</type>
<position>-42,-214</position>
<input>
<ID>IN_0</ID>852 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add12</lparam></gate>
<gate>
<ID>505</ID>
<type>DA_FROM</type>
<position>-42,-152.5</position>
<input>
<ID>IN_0</ID>654 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>543</ID>
<type>AA_AND2</type>
<position>-36,-188.5</position>
<input>
<ID>IN_0</ID>678 </input>
<input>
<ID>IN_1</ID>685 </input>
<output>
<ID>OUT</ID>677 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>506</ID>
<type>DA_FROM</type>
<position>-42,-157.5</position>
<input>
<ID>IN_0</ID>655 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>507</ID>
<type>AA_AND2</type>
<position>-36,-158.5</position>
<input>
<ID>IN_0</ID>655 </input>
<input>
<ID>IN_1</ID>657 </input>
<output>
<ID>OUT</ID>656 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>685</ID>
<type>DA_FROM</type>
<position>13,-212</position>
<input>
<ID>IN_0</ID>825 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>508</ID>
<type>DA_FROM</type>
<position>-42,-159.5</position>
<input>
<ID>IN_0</ID>657 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID InpR4</lparam></gate>
<gate>
<ID>716</ID>
<type>AE_SMALL_INVERTER</type>
<position>-51,-224</position>
<input>
<ID>IN_0</ID>849 </input>
<output>
<ID>OUT_0</ID>857 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>509</ID>
<type>DA_FROM</type>
<position>-42,-149.5</position>
<input>
<ID>IN_0</ID>659 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo5</lparam></gate>
<gate>
<ID>531</ID>
<type>AA_AND2</type>
<position>-50,-169.5</position>
<input>
<ID>IN_0</ID>666 </input>
<input>
<ID>IN_1</ID>667 </input>
<output>
<ID>OUT</ID>664 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>510</ID>
<type>DA_FROM</type>
<position>-42,-154.5</position>
<input>
<ID>IN_0</ID>660 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo3</lparam></gate>
<gate>
<ID>514</ID>
<type>AA_AND2</type>
<position>74,-168.5</position>
<input>
<ID>IN_0</ID>717 </input>
<input>
<ID>IN_1</ID>716 </input>
<output>
<ID>OUT</ID>715 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>516</ID>
<type>DA_FROM</type>
<position>-3,-208</position>
<input>
<ID>IN_0</ID>822 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR13</lparam></gate>
<gate>
<ID>518</ID>
<type>FF_GND</type>
<position>-27.5,-179.5</position>
<output>
<ID>OUT_0</ID>684 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>520</ID>
<type>DA_FROM</type>
<position>68,-167.5</position>
<input>
<ID>IN_0</ID>717 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>524</ID>
<type>AA_AND2</type>
<position>74,-178.5</position>
<input>
<ID>IN_0</ID>725 </input>
<input>
<ID>IN_1</ID>718 </input>
<output>
<ID>OUT</ID>724 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>528</ID>
<type>DE_TO</type>
<position>-16.5,-183.5</position>
<input>
<ID>IN_0</ID>668 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi8</lparam></gate>
<gate>
<ID>532</ID>
<type>DA_FROM</type>
<position>-42,-167.5</position>
<input>
<ID>IN_0</ID>665 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>536</ID>
<type>DA_FROM</type>
<position>-42,-172.5</position>
<input>
<ID>IN_0</ID>669 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>540</ID>
<type>AA_AND2</type>
<position>-36,-183.5</position>
<input>
<ID>IN_0</ID>676 </input>
<input>
<ID>IN_1</ID>675 </input>
<output>
<ID>OUT</ID>674 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>544</ID>
<type>DA_FROM</type>
<position>-42,-187.5</position>
<input>
<ID>IN_0</ID>678 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>556</ID>
<type>DE_OR8</type>
<position>31.5,-183.5</position>
<input>
<ID>IN_0</ID>710 </input>
<input>
<ID>IN_1</ID>689 </input>
<input>
<ID>IN_2</ID>697 </input>
<input>
<ID>IN_3</ID>698 </input>
<input>
<ID>IN_4</ID>872 </input>
<input>
<ID>IN_5</ID>705 </input>
<input>
<ID>IN_6</ID>703 </input>
<input>
<ID>IN_7</ID>700 </input>
<output>
<ID>OUT</ID>694 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>558</ID>
<type>AA_AND2</type>
<position>5,-169.5</position>
<input>
<ID>IN_0</ID>692 </input>
<input>
<ID>IN_1</ID>693 </input>
<output>
<ID>OUT</ID>690 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>560</ID>
<type>DA_FROM</type>
<position>-3,-168.5</position>
<input>
<ID>IN_0</ID>692 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR9</lparam></gate>
<gate>
<ID>562</ID>
<type>AA_AND2</type>
<position>19,-173.5</position>
<input>
<ID>IN_0</ID>695 </input>
<input>
<ID>IN_1</ID>696 </input>
<output>
<ID>OUT</ID>697 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>564</ID>
<type>DA_FROM</type>
<position>13,-174.5</position>
<input>
<ID>IN_0</ID>696 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add9</lparam></gate>
<gate>
<ID>566</ID>
<type>DA_FROM</type>
<position>13,-177.5</position>
<input>
<ID>IN_0</ID>699 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>568</ID>
<type>AE_SMALL_INVERTER</type>
<position>4,-184.5</position>
<input>
<ID>IN_0</ID>693 </input>
<output>
<ID>OUT_0</ID>701 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>572</ID>
<type>AA_AND2</type>
<position>19,-193.5</position>
<input>
<ID>IN_0</ID>706 </input>
<input>
<ID>IN_1</ID>712 </input>
<output>
<ID>OUT</ID>705 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>578</ID>
<type>FF_GND</type>
<position>82.5,-179.5</position>
<output>
<ID>OUT_0</ID>736 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>579</ID>
<type>DE_OR8</type>
<position>86.5,-183.5</position>
<input>
<ID>IN_0</ID>736 </input>
<input>
<ID>IN_1</ID>715 </input>
<input>
<ID>IN_2</ID>723 </input>
<input>
<ID>IN_3</ID>724 </input>
<input>
<ID>IN_4</ID>873 </input>
<input>
<ID>IN_5</ID>731 </input>
<input>
<ID>IN_6</ID>729 </input>
<input>
<ID>IN_7</ID>726 </input>
<output>
<ID>OUT</ID>720 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>582</ID>
<type>DA_FROM</type>
<position>52,-170.5</position>
<input>
<ID>IN_0</ID>719 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo10</lparam></gate>
<gate>
<ID>583</ID>
<type>AA_AND2</type>
<position>74,-173.5</position>
<input>
<ID>IN_0</ID>721 </input>
<input>
<ID>IN_1</ID>722 </input>
<output>
<ID>OUT</ID>723 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>586</ID>
<type>AE_SMALL_INVERTER</type>
<position>59,-184.5</position>
<input>
<ID>IN_0</ID>719 </input>
<output>
<ID>OUT_0</ID>727 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>587</ID>
<type>AA_AND2</type>
<position>74,-188.5</position>
<input>
<ID>IN_0</ID>730 </input>
<input>
<ID>IN_1</ID>737 </input>
<output>
<ID>OUT</ID>729 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>590</ID>
<type>DA_FROM</type>
<position>68,-192.5</position>
<input>
<ID>IN_0</ID>732 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>594</ID>
<type>DA_FROM</type>
<position>68,-194.5</position>
<input>
<ID>IN_0</ID>738 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo9</lparam></gate>
<gate>
<ID>598</ID>
<type>DE_TO</type>
<position>148.5,-183.5</position>
<input>
<ID>IN_0</ID>746 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi11</lparam></gate>
<gate>
<ID>599</ID>
<type>DE_OR8</type>
<position>141.5,-183.5</position>
<input>
<ID>IN_0</ID>762 </input>
<input>
<ID>IN_1</ID>741 </input>
<input>
<ID>IN_2</ID>749 </input>
<input>
<ID>IN_3</ID>750 </input>
<input>
<ID>IN_4</ID>874 </input>
<input>
<ID>IN_5</ID>757 </input>
<input>
<ID>IN_6</ID>755 </input>
<input>
<ID>IN_7</ID>752 </input>
<output>
<ID>OUT</ID>746 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>600</ID>
<type>AA_AND2</type>
<position>129,-168.5</position>
<input>
<ID>IN_0</ID>743 </input>
<input>
<ID>IN_1</ID>742 </input>
<output>
<ID>OUT</ID>741 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>602</ID>
<type>DA_FROM</type>
<position>123,-167.5</position>
<input>
<ID>IN_0</ID>743 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>604</ID>
<type>DA_FROM</type>
<position>107,-170.5</position>
<input>
<ID>IN_0</ID>745 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo11</lparam></gate>
<gate>
<ID>606</ID>
<type>DA_FROM</type>
<position>123,-172.5</position>
<input>
<ID>IN_0</ID>747 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>607</ID>
<type>DA_FROM</type>
<position>123,-174.5</position>
<input>
<ID>IN_0</ID>748 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add11</lparam></gate>
<gate>
<ID>608</ID>
<type>AA_AND2</type>
<position>129,-178.5</position>
<input>
<ID>IN_0</ID>751 </input>
<input>
<ID>IN_1</ID>744 </input>
<output>
<ID>OUT</ID>750 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>610</ID>
<type>AA_AND2</type>
<position>129,-183.5</position>
<input>
<ID>IN_0</ID>754 </input>
<input>
<ID>IN_1</ID>753 </input>
<output>
<ID>OUT</ID>752 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>612</ID>
<type>DA_FROM</type>
<position>123,-182.5</position>
<input>
<ID>IN_0</ID>754 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>614</ID>
<type>DA_FROM</type>
<position>123,-187.5</position>
<input>
<ID>IN_0</ID>756 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>616</ID>
<type>DA_FROM</type>
<position>123,-192.5</position>
<input>
<ID>IN_0</ID>758 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>620</ID>
<type>DA_FROM</type>
<position>123,-189.5</position>
<input>
<ID>IN_0</ID>763 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo12</lparam></gate>
<gate>
<ID>624</ID>
<type>FF_GND</type>
<position>137.5,-219</position>
<output>
<ID>OUT_0</ID>788 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>626</ID>
<type>DE_OR8</type>
<position>141.5,-223</position>
<input>
<ID>IN_0</ID>788 </input>
<input>
<ID>IN_1</ID>767 </input>
<input>
<ID>IN_2</ID>775 </input>
<input>
<ID>IN_3</ID>776 </input>
<input>
<ID>IN_4</ID>878 </input>
<input>
<ID>IN_5</ID>783 </input>
<input>
<ID>IN_6</ID>781 </input>
<input>
<ID>IN_7</ID>778 </input>
<output>
<ID>OUT</ID>772 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>628</ID>
<type>AA_AND2</type>
<position>115,-209</position>
<input>
<ID>IN_0</ID>770 </input>
<input>
<ID>IN_1</ID>771 </input>
<output>
<ID>OUT</ID>768 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>630</ID>
<type>DA_FROM</type>
<position>107,-208</position>
<input>
<ID>IN_0</ID>770 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR15</lparam></gate>
<gate>
<ID>632</ID>
<type>AA_AND2</type>
<position>129,-213</position>
<input>
<ID>IN_0</ID>773 </input>
<input>
<ID>IN_1</ID>774 </input>
<output>
<ID>OUT</ID>775 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>634</ID>
<type>DA_FROM</type>
<position>123,-214</position>
<input>
<ID>IN_0</ID>774 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add15</lparam></gate>
<gate>
<ID>636</ID>
<type>DA_FROM</type>
<position>123,-217</position>
<input>
<ID>IN_0</ID>777 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>638</ID>
<type>AE_SMALL_INVERTER</type>
<position>114,-224</position>
<input>
<ID>IN_0</ID>771 </input>
<output>
<ID>OUT_0</ID>779 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>642</ID>
<type>AA_AND2</type>
<position>129,-233</position>
<input>
<ID>IN_0</ID>784 </input>
<input>
<ID>IN_1</ID>790 </input>
<output>
<ID>OUT</ID>783 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>643</ID>
<type>DA_FROM</type>
<position>123,-232</position>
<input>
<ID>IN_0</ID>784 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>647</ID>
<type>DA_FROM</type>
<position>123,-229</position>
<input>
<ID>IN_0</ID>789 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>651</ID>
<type>FF_GND</type>
<position>82.5,-219</position>
<output>
<ID>OUT_0</ID>814 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>654</ID>
<type>AA_AND2</type>
<position>74,-208</position>
<input>
<ID>IN_0</ID>795 </input>
<input>
<ID>IN_1</ID>794 </input>
<output>
<ID>OUT</ID>793 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>655</ID>
<type>AA_AND2</type>
<position>60,-209</position>
<input>
<ID>IN_0</ID>796 </input>
<input>
<ID>IN_1</ID>797 </input>
<output>
<ID>OUT</ID>794 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>656</ID>
<type>DA_FROM</type>
<position>68,-207</position>
<input>
<ID>IN_0</ID>795 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>658</ID>
<type>DA_FROM</type>
<position>52,-210</position>
<input>
<ID>IN_0</ID>797 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo14</lparam></gate>
<gate>
<ID>659</ID>
<type>AA_AND2</type>
<position>74,-213</position>
<input>
<ID>IN_0</ID>799 </input>
<input>
<ID>IN_1</ID>800 </input>
<output>
<ID>OUT</ID>801 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>662</ID>
<type>AA_AND2</type>
<position>74,-218</position>
<input>
<ID>IN_0</ID>803 </input>
<input>
<ID>IN_1</ID>796 </input>
<output>
<ID>OUT</ID>802 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>663</ID>
<type>DA_FROM</type>
<position>68,-217</position>
<input>
<ID>IN_0</ID>803 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>666</ID>
<type>DA_FROM</type>
<position>68,-222</position>
<input>
<ID>IN_0</ID>806 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>667</ID>
<type>AA_AND2</type>
<position>74,-228</position>
<input>
<ID>IN_0</ID>808 </input>
<input>
<ID>IN_1</ID>815 </input>
<output>
<ID>OUT</ID>807 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>674</ID>
<type>DA_FROM</type>
<position>68,-234</position>
<input>
<ID>IN_0</ID>816 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo13</lparam></gate>
<gate>
<ID>678</ID>
<type>DE_TO</type>
<position>38.5,-223</position>
<input>
<ID>IN_0</ID>824 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi13</lparam></gate>
<gate>
<ID>679</ID>
<type>DE_OR8</type>
<position>31.5,-223</position>
<input>
<ID>IN_0</ID>840 </input>
<input>
<ID>IN_1</ID>819 </input>
<input>
<ID>IN_2</ID>827 </input>
<input>
<ID>IN_3</ID>828 </input>
<input>
<ID>IN_4</ID>876 </input>
<input>
<ID>IN_5</ID>835 </input>
<input>
<ID>IN_6</ID>833 </input>
<input>
<ID>IN_7</ID>830 </input>
<output>
<ID>OUT</ID>824 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>682</ID>
<type>DA_FROM</type>
<position>13,-207</position>
<input>
<ID>IN_0</ID>821 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>683</ID>
<type>DA_FROM</type>
<position>-3,-210</position>
<input>
<ID>IN_0</ID>823 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo13</lparam></gate>
<gate>
<ID>686</ID>
<type>DA_FROM</type>
<position>13,-214</position>
<input>
<ID>IN_0</ID>826 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID add13</lparam></gate>
<gate>
<ID>687</ID>
<type>AA_AND2</type>
<position>19,-218</position>
<input>
<ID>IN_0</ID>829 </input>
<input>
<ID>IN_1</ID>822 </input>
<output>
<ID>OUT</ID>828 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>690</ID>
<type>AE_SMALL_INVERTER</type>
<position>4,-224</position>
<input>
<ID>IN_0</ID>823 </input>
<output>
<ID>OUT_0</ID>831 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>691</ID>
<type>DA_FROM</type>
<position>13,-222</position>
<input>
<ID>IN_0</ID>832 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>694</ID>
<type>AA_AND2</type>
<position>19,-233</position>
<input>
<ID>IN_0</ID>836 </input>
<input>
<ID>IN_1</ID>842 </input>
<output>
<ID>OUT</ID>835 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>695</ID>
<type>DA_FROM</type>
<position>13,-232</position>
<input>
<ID>IN_0</ID>836 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>699</ID>
<type>DA_FROM</type>
<position>13,-229</position>
<input>
<ID>IN_0</ID>841 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo14</lparam></gate>
<gate>
<ID>702</ID>
<type>FF_GND</type>
<position>-27.5,-219</position>
<output>
<ID>OUT_0</ID>866 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>703</ID>
<type>DE_TO</type>
<position>-16.5,-223</position>
<input>
<ID>IN_0</ID>850 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACi12</lparam></gate>
<gate>
<ID>705</ID>
<type>AA_AND2</type>
<position>-36,-208</position>
<input>
<ID>IN_0</ID>847 </input>
<input>
<ID>IN_1</ID>846 </input>
<output>
<ID>OUT</ID>845 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>707</ID>
<type>DA_FROM</type>
<position>-42,-207</position>
<input>
<ID>IN_0</ID>847 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>709</ID>
<type>DA_FROM</type>
<position>-58,-210</position>
<input>
<ID>IN_0</ID>849 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo12</lparam></gate>
<gate>
<ID>713</ID>
<type>AA_AND2</type>
<position>-36,-218</position>
<input>
<ID>IN_0</ID>855 </input>
<input>
<ID>IN_1</ID>848 </input>
<output>
<ID>OUT</ID>854 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>715</ID>
<type>AA_AND2</type>
<position>-36,-223</position>
<input>
<ID>IN_0</ID>858 </input>
<input>
<ID>IN_1</ID>857 </input>
<output>
<ID>OUT</ID>856 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>717</ID>
<type>DA_FROM</type>
<position>-42,-222</position>
<input>
<ID>IN_0</ID>858 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>719</ID>
<type>DA_FROM</type>
<position>-42,-227</position>
<input>
<ID>IN_0</ID>860 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>721</ID>
<type>DA_FROM</type>
<position>-42,-232</position>
<input>
<ID>IN_0</ID>862 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>725</ID>
<type>DA_FROM</type>
<position>-42,-229</position>
<input>
<ID>IN_0</ID>867 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo13</lparam></gate>
<gate>
<ID>738</ID>
<type>FF_GND</type>
<position>-27.5,-228.5</position>
<output>
<ID>OUT_0</ID>875 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1047</ID>
<type>AE_SMALL_INVERTER</type>
<position>-100,-161</position>
<input>
<ID>IN_0</ID>348 </input>
<output>
<ID>OUT_0</ID>1177 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>-103.5,-164.5</position>
<gparam>LABEL_TEXT ALU</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>266 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-127,-105,-127</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>746 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145.5,-183.5,146.5,-183.5</points>
<connection>
<GID>599</GID>
<name>OUT</name></connection>
<connection>
<GID>598</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-128,-105,-128</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>538 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-127.5,71,-127.5</points>
<connection>
<GID>437</GID>
<name>IN_0</name></connection>
<connection>
<GID>435</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>208 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102,-141,-102,-140</points>
<connection>
<GID>156</GID>
<name>carry_out</name></connection>
<connection>
<GID>157</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>447 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-88,71,-88</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<connection>
<GID>354</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>738 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-194.5,71,-194.5</points>
<connection>
<GID>589</GID>
<name>IN_1</name></connection>
<connection>
<GID>594</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-144,-105,-144</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_B_0</name></connection></hsegment></shape></wire>
<wire>
<ID>318 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-137,-105,-137</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>446 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-90,71,-90</points>
<connection>
<GID>355</GID>
<name>OUT</name></connection>
<connection>
<GID>354</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-97.5,-86.5,-97.5</points>
<connection>
<GID>154</GID>
<name>OUT_1</name></connection>
<connection>
<GID>162</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>628 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-152.5,16,-152.5</points>
<connection>
<GID>478</GID>
<name>IN_0</name></connection>
<connection>
<GID>477</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-100,-105,-100</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<connection>
<GID>206</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>851 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-212,-39,-212</points>
<connection>
<GID>711</GID>
<name>IN_0</name></connection>
<connection>
<GID>710</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>652 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-147.5,-39,-147.5</points>
<connection>
<GID>503</GID>
<name>IN_0</name></connection>
<connection>
<GID>502</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>445 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-101.5,81,-89</points>
<intersection>-101.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-89,81,-89</points>
<connection>
<GID>354</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-101.5,83.5,-101.5</points>
<connection>
<GID>353</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>251 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-114.5,-86.5,-114.5</points>
<connection>
<GID>177</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>758 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-192.5,126,-192.5</points>
<connection>
<GID>615</GID>
<name>IN_0</name></connection>
<connection>
<GID>616</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-94,-105,-94</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<connection>
<GID>154</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>614 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-128.5,2,-128.5</points>
<connection>
<GID>463</GID>
<name>IN_0</name></connection>
<connection>
<GID>465</GID>
<name>IN_0</name></connection>
<intersection>1 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1,-139.5,1,-128.5</points>
<intersection>-139.5 8</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>1,-139.5,16,-139.5</points>
<connection>
<GID>470</GID>
<name>IN_1</name></connection>
<intersection>1 7</intersection></hsegment></shape></wire>
<wire>
<ID>608 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-154.5,71,-154.5</points>
<connection>
<GID>450</GID>
<name>IN_1</name></connection>
<connection>
<GID>456</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-111,-105,-111</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>IN_B_1</name></connection></hsegment></shape></wire>
<wire>
<ID>600 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-147.5,71,-147.5</points>
<connection>
<GID>449</GID>
<name>IN_0</name></connection>
<connection>
<GID>448</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-129,-105,-129</points>
<connection>
<GID>156</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>199</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>329 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-89,-53,-89</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>-54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-54,-100,-54,-89</points>
<intersection>-100 8</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-54,-100,-39,-100</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>-54 7</intersection></hsegment></shape></wire>
<wire>
<ID>664 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-169.5,-39,-169.5</points>
<connection>
<GID>530</GID>
<name>IN_1</name></connection>
<connection>
<GID>531</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>728 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-182.5,71,-182.5</points>
<connection>
<GID>522</GID>
<name>IN_0</name></connection>
<connection>
<GID>526</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>301 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-101,-105,-101</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-102,-105,-102</points>
<connection>
<GID>154</GID>
<name>IN_2</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>302 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-103,-105,-103</points>
<connection>
<GID>154</GID>
<name>IN_3</name></connection>
<connection>
<GID>209</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-93,-105,-93</points>
<connection>
<GID>154</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>828 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-222.5,25,-218</points>
<intersection>-222.5 1</intersection>
<intersection>-218 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-222.5,28.5,-222.5</points>
<connection>
<GID>679</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-218,25,-218</points>
<connection>
<GID>687</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>667 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-170.5,-53,-170.5</points>
<connection>
<GID>531</GID>
<name>IN_1</name></connection>
<connection>
<GID>534</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-55,-184.5,-55,-170.5</points>
<intersection>-184.5 6</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-55,-184.5,-53,-184.5</points>
<connection>
<GID>541</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-95,-105,-95</points>
<connection>
<GID>154</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>191</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-96,-105,-96</points>
<connection>
<GID>154</GID>
<name>IN_B_3</name></connection>
<connection>
<GID>192</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>298 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-134,-105,-134</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>209 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102,-90,-102,-87</points>
<connection>
<GID>154</GID>
<name>carry_in</name></connection>
<intersection>-87 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>-100.5,-88,-100.5,-87</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-87 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-102,-87,-100.5,-87</points>
<intersection>-102 0</intersection>
<intersection>-100.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>245 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-96.5,-96,-96.5</points>
<connection>
<GID>154</GID>
<name>OUT_0</name></connection>
<connection>
<GID>161</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>270 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-147,-105,-147</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>779 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-224,126,-224</points>
<connection>
<GID>637</GID>
<name>IN_1</name></connection>
<connection>
<GID>638</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>246 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-98.5,-96,-98.5</points>
<connection>
<GID>154</GID>
<name>OUT_2</name></connection>
<connection>
<GID>164</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>253 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-99.5,-86.5,-99.5</points>
<connection>
<GID>154</GID>
<name>OUT_3</name></connection>
<connection>
<GID>166</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>867 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-229,-39,-229</points>
<connection>
<GID>718</GID>
<name>IN_1</name></connection>
<connection>
<GID>725</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>206 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102,-107,-102,-106</points>
<connection>
<GID>154</GID>
<name>carry_out</name></connection>
<connection>
<GID>155</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>808 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-227,71,-227</points>
<connection>
<GID>517</GID>
<name>IN_0</name></connection>
<connection>
<GID>667</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>663 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-181,-29,-168.5</points>
<intersection>-181 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,-168.5,-29,-168.5</points>
<connection>
<GID>530</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29,-181,-26.5,-181</points>
<connection>
<GID>529</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>872 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-188,27.5,-187</points>
<connection>
<GID>732</GID>
<name>OUT_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-187,28.5,-187</points>
<connection>
<GID>556</GID>
<name>IN_4</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>727 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-184.5,71,-184.5</points>
<connection>
<GID>522</GID>
<name>IN_1</name></connection>
<connection>
<GID>586</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>299 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-120,-105,-120</points>
<connection>
<GID>155</GID>
<name>IN_3</name></connection>
<connection>
<GID>213</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>726 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-184,80,-183.5</points>
<intersection>-184 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-184,83.5,-184</points>
<connection>
<GID>579</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-183.5,80,-183.5</points>
<connection>
<GID>522</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-113,-105,-113</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<connection>
<GID>155</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>296 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-151,-105,-151</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>665 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-167.5,-39,-167.5</points>
<connection>
<GID>530</GID>
<name>IN_0</name></connection>
<connection>
<GID>532</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-150.5,-86.5,-150.5</points>
<connection>
<GID>157</GID>
<name>OUT_3</name></connection>
<connection>
<GID>187</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-130,-105,-130</points>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_B_3</name></connection></hsegment></shape></wire>
<wire>
<ID>414 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-100.5,-26.5,-98.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-98.5,-26.5,-98.5</points>
<intersection>-27.5 3</intersection>
<intersection>-26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-99,-27.5,-98.5</points>
<connection>
<GID>316</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>654 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-152.5,-39,-152.5</points>
<connection>
<GID>505</GID>
<name>IN_0</name></connection>
<connection>
<GID>504</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-117,-105,-117</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>300 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-118,-105,-118</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<connection>
<GID>211</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-119,-105,-119</points>
<connection>
<GID>155</GID>
<name>IN_2</name></connection>
<connection>
<GID>212</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>750 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-183,135,-178.5</points>
<intersection>-183 1</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-183,138.5,-183</points>
<connection>
<GID>599</GID>
<name>IN_3</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-178.5,135,-178.5</points>
<connection>
<GID>608</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-110,-105,-110</points>
<connection>
<GID>155</GID>
<name>IN_B_0</name></connection>
<connection>
<GID>193</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-112,-105,-112</points>
<connection>
<GID>155</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>195</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>244 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-113.5,-96,-113.5</points>
<connection>
<GID>155</GID>
<name>OUT_0</name></connection>
<connection>
<GID>176</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-115.5,-96,-115.5</points>
<connection>
<GID>155</GID>
<name>OUT_2</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>252 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-116.5,-86.5,-116.5</points>
<connection>
<GID>155</GID>
<name>OUT_3</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>529 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-158.5,136,-147</points>
<intersection>-158.5 2</intersection>
<intersection>-147 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-147,138.5,-147</points>
<connection>
<GID>407</GID>
<name>IN_4</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-158.5,136,-158.5</points>
<connection>
<GID>426</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>207 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102,-124,-102,-123</points>
<connection>
<GID>155</GID>
<name>carry_out</name></connection>
<connection>
<GID>156</GID>
<name>carry_in</name></connection></vsegment></shape></wire>
<wire>
<ID>512 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-144,135,-143.5</points>
<intersection>-144 1</intersection>
<intersection>-143.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-144,138.5,-144</points>
<connection>
<GID>407</GID>
<name>IN_7</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-143.5,135,-143.5</points>
<connection>
<GID>418</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>305 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-135,-105,-135</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<connection>
<GID>215</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>632 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-140,28.5,-138</points>
<connection>
<GID>461</GID>
<name>IN_0</name></connection>
<intersection>-138 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-138,28.5,-138</points>
<intersection>27.5 3</intersection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-138.5,27.5,-138</points>
<connection>
<GID>459</GID>
<name>OUT_0</name></connection>
<intersection>-138 2</intersection></vsegment></shape></wire>
<wire>
<ID>297 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-136,-105,-136</points>
<connection>
<GID>156</GID>
<name>IN_2</name></connection>
<connection>
<GID>216</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>247 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-130.5,-96,-130.5</points>
<connection>
<GID>156</GID>
<name>OUT_0</name></connection>
<connection>
<GID>180</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-146,-105,-146</points>
<connection>
<GID>157</GID>
<name>IN_B_2</name></connection>
<connection>
<GID>203</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-131.5,-86.5,-131.5</points>
<connection>
<GID>156</GID>
<name>OUT_1</name></connection>
<connection>
<GID>181</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>642 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-143.5,-18.5,-143.5</points>
<connection>
<GID>488</GID>
<name>OUT</name></connection>
<connection>
<GID>487</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-106,-153,-105,-153</points>
<connection>
<GID>157</GID>
<name>IN_2</name></connection>
<connection>
<GID>224</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>248 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-132.5,-96,-132.5</points>
<connection>
<GID>156</GID>
<name>OUT_2</name></connection>
<connection>
<GID>182</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-133.5,-86.5,-133.5</points>
<connection>
<GID>156</GID>
<name>OUT_3</name></connection>
<connection>
<GID>183</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>508 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-134.5,126,-134.5</points>
<connection>
<GID>413</GID>
<name>IN_1</name></connection>
<connection>
<GID>415</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>685 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-189.5,-39,-189.5</points>
<connection>
<GID>543</GID>
<name>IN_1</name></connection>
<connection>
<GID>550</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>304 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-152,-105,-152</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<connection>
<GID>222</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>650 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-142.5,-39,-142.5</points>
<connection>
<GID>501</GID>
<name>IN_0</name></connection>
<connection>
<GID>499</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>303 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-115.5,-154,-105,-154</points>
<connection>
<GID>157</GID>
<name>IN_3</name></connection>
<connection>
<GID>226</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>604 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-158.5,81,-147</points>
<intersection>-158.5 2</intersection>
<intersection>-147 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-147,83.5,-147</points>
<connection>
<GID>434</GID>
<name>IN_4</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-158.5,81,-158.5</points>
<connection>
<GID>453</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-114,-145,-105,-145</points>
<connection>
<GID>157</GID>
<name>IN_B_1</name></connection>
<connection>
<GID>202</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>249 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-147.5,-96,-147.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-148.5,-86.5,-148.5</points>
<connection>
<GID>157</GID>
<name>OUT_1</name></connection>
<connection>
<GID>185</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>799 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-212,71,-212</points>
<connection>
<GID>660</GID>
<name>IN_0</name></connection>
<connection>
<GID>659</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>250 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-97,-149.5,-96,-149.5</points>
<connection>
<GID>157</GID>
<name>OUT_2</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>525 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-147.5,126,-147.5</points>
<connection>
<GID>422</GID>
<name>IN_0</name></connection>
<connection>
<GID>421</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>348 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-102,-161,-102,-157</points>
<connection>
<GID>1047</GID>
<name>IN_0</name></connection>
<connection>
<GID>157</GID>
<name>carry_out</name></connection>
<intersection>-158.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-102,-158.5,-97,-158.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>-102 0</intersection></hsegment></shape></wire>
<wire>
<ID>334 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-102.5,-29.5,-94</points>
<intersection>-102.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-102.5,-26.5,-102.5</points>
<connection>
<GID>233</GID>
<name>IN_2</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-94,-29.5,-94</points>
<connection>
<GID>260</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-98,-161,-97,-161</points>
<connection>
<GID>1047</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1048</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>439 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-120,16,-120</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<connection>
<GID>346</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>666 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-168.5,-53,-168.5</points>
<connection>
<GID>531</GID>
<name>IN_0</name></connection>
<connection>
<GID>533</GID>
<name>IN_0</name></connection>
<intersection>-54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-54,-179.5,-54,-168.5</points>
<intersection>-179.5 8</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-54,-179.5,-39,-179.5</points>
<connection>
<GID>538</GID>
<name>IN_1</name></connection>
<intersection>-54 7</intersection></hsegment></shape></wire>
<wire>
<ID>644 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-134.5,-39,-134.5</points>
<connection>
<GID>494</GID>
<name>IN_1</name></connection>
<connection>
<GID>496</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>437 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-118,16,-118</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<connection>
<GID>344</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>675 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-184.5,-39,-184.5</points>
<connection>
<GID>541</GID>
<name>OUT_0</name></connection>
<connection>
<GID>540</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>623 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-144.5,16,-144.5</points>
<connection>
<GID>473</GID>
<name>OUT_0</name></connection>
<connection>
<GID>472</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>458 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-103,71,-103</points>
<connection>
<GID>366</GID>
<name>IN_0</name></connection>
<connection>
<GID>364</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>457 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-105,71,-105</points>
<connection>
<GID>365</GID>
<name>OUT_0</name></connection>
<connection>
<GID>364</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>456 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-104.5,80,-104</points>
<intersection>-104.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-104.5,83.5,-104.5</points>
<connection>
<GID>353</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-104,80,-104</points>
<connection>
<GID>364</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>684 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-180,-26.5,-178</points>
<connection>
<GID>529</GID>
<name>IN_0</name></connection>
<intersection>-178 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-178,-26.5,-178</points>
<intersection>-27.5 3</intersection>
<intersection>-26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-178.5,-27.5,-178</points>
<connection>
<GID>518</GID>
<name>OUT_0</name></connection>
<intersection>-178 2</intersection></vsegment></shape></wire>
<wire>
<ID>816 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-234,71,-234</points>
<connection>
<GID>668</GID>
<name>IN_1</name></connection>
<connection>
<GID>674</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>671 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-182,-29.5,-173.5</points>
<intersection>-182 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-182,-26.5,-182</points>
<connection>
<GID>529</GID>
<name>IN_2</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-173.5,-29.5,-173.5</points>
<connection>
<GID>535</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>672 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-183,-30,-178.5</points>
<intersection>-183 1</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-183,-26.5,-183</points>
<connection>
<GID>529</GID>
<name>IN_3</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-178.5,-30,-178.5</points>
<connection>
<GID>538</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>871 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-188,-27.5,-187</points>
<connection>
<GID>730</GID>
<name>OUT_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,-187,-26.5,-187</points>
<connection>
<GID>529</GID>
<name>IN_4</name></connection>
<intersection>-27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>824 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-223,36.5,-223</points>
<connection>
<GID>679</GID>
<name>OUT</name></connection>
<connection>
<GID>678</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>679 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-193.5,-29.5,-186</points>
<intersection>-193.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-186,-26.5,-186</points>
<connection>
<GID>529</GID>
<name>IN_5</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-193.5,-29.5,-193.5</points>
<connection>
<GID>545</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>830 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-223.5,25,-223</points>
<intersection>-223.5 1</intersection>
<intersection>-223 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-223.5,28.5,-223.5</points>
<connection>
<GID>679</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-223,25,-223</points>
<connection>
<GID>689</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>677 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-188.5,-30,-185</points>
<intersection>-188.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-185,-26.5,-185</points>
<connection>
<GID>529</GID>
<name>IN_6</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-188.5,-30,-188.5</points>
<connection>
<GID>543</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>674 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-184,-30,-183.5</points>
<intersection>-184 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-184,-26.5,-184</points>
<connection>
<GID>529</GID>
<name>IN_7</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-183.5,-30,-183.5</points>
<connection>
<GID>540</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>333 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-95,-39,-95</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<connection>
<GID>260</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>668 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-183.5,-18.5,-183.5</points>
<connection>
<GID>529</GID>
<name>OUT</name></connection>
<connection>
<GID>528</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>615 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-130.5,2,-130.5</points>
<connection>
<GID>463</GID>
<name>IN_1</name></connection>
<connection>
<GID>466</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>0,-144.5,0,-130.5</points>
<intersection>-144.5 6</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>0,-144.5,2,-144.5</points>
<connection>
<GID>473</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment></shape></wire>
<wire>
<ID>450 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-104,91.5,-104</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<connection>
<GID>352</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>496 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-100.5,138.5,-98.5</points>
<connection>
<GID>380</GID>
<name>IN_0</name></connection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-98.5,138.5,-98.5</points>
<intersection>137.5 3</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>137.5,-99,137.5,-98.5</points>
<connection>
<GID>378</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>826 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-214,16,-214</points>
<connection>
<GID>684</GID>
<name>IN_1</name></connection>
<connection>
<GID>686</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>673 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-177.5,-39,-177.5</points>
<connection>
<GID>538</GID>
<name>IN_0</name></connection>
<connection>
<GID>539</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>777 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-217,126,-217</points>
<connection>
<GID>635</GID>
<name>IN_0</name></connection>
<connection>
<GID>636</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>455 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-98,71,-98</points>
<connection>
<GID>363</GID>
<name>IN_0</name></connection>
<connection>
<GID>362</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>753 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-184.5,126,-184.5</points>
<connection>
<GID>611</GID>
<name>OUT_0</name></connection>
<connection>
<GID>610</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>778 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-223.5,135,-223</points>
<intersection>-223.5 1</intersection>
<intersection>-223 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-223.5,138.5,-223.5</points>
<connection>
<GID>626</GID>
<name>IN_7</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-223,135,-223</points>
<connection>
<GID>637</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>448 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-89,57,-89</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>56,-100,56,-89</points>
<intersection>-100 8</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>56,-100,71,-100</points>
<connection>
<GID>362</GID>
<name>IN_1</name></connection>
<intersection>56 7</intersection></hsegment></shape></wire>
<wire>
<ID>603 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-157.5,71,-157.5</points>
<connection>
<GID>452</GID>
<name>IN_0</name></connection>
<connection>
<GID>453</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>454 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-103.5,80,-99</points>
<intersection>-103.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-103.5,83.5,-103.5</points>
<connection>
<GID>353</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-99,80,-99</points>
<connection>
<GID>362</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>463 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-118,71,-118</points>
<connection>
<GID>371</GID>
<name>IN_0</name></connection>
<connection>
<GID>372</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>465 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-120,71,-120</points>
<connection>
<GID>372</GID>
<name>IN_1</name></connection>
<connection>
<GID>373</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>794 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-209,71,-209</points>
<connection>
<GID>654</GID>
<name>IN_1</name></connection>
<connection>
<GID>655</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>641 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-130.5,-53,-130.5</points>
<connection>
<GID>490</GID>
<name>IN_1</name></connection>
<connection>
<GID>493</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-55,-144.5,-55,-130.5</points>
<intersection>-144.5 6</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-55,-144.5,-53,-144.5</points>
<connection>
<GID>500</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment></shape></wire>
<wire>
<ID>464 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-119,81,-107.5</points>
<intersection>-119 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81,-107.5,83.5,-107.5</points>
<connection>
<GID>353</GID>
<name>IN_4</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-119,81,-119</points>
<connection>
<GID>372</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>341 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-109,-30,-105.5</points>
<intersection>-109 2</intersection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-105.5,-26.5,-105.5</points>
<connection>
<GID>233</GID>
<name>IN_6</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-109,-30,-109</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>676 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-182.5,-39,-182.5</points>
<connection>
<GID>542</GID>
<name>IN_0</name></connection>
<connection>
<GID>540</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>789 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-229,126,-229</points>
<connection>
<GID>640</GID>
<name>IN_1</name></connection>
<connection>
<GID>647</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>451 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-93,71,-93</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<connection>
<GID>360</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>670 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-174.5,-39,-174.5</points>
<connection>
<GID>535</GID>
<name>IN_1</name></connection>
<connection>
<GID>537</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>345 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-118,-39,-118</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<connection>
<GID>286</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>680 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-192.5,-39,-192.5</points>
<connection>
<GID>546</GID>
<name>IN_0</name></connection>
<connection>
<GID>545</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>347 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-120,-39,-120</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<connection>
<GID>290</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>710 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-180,28.5,-178</points>
<connection>
<GID>556</GID>
<name>IN_0</name></connection>
<intersection>-178 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-178,28.5,-178</points>
<intersection>27.5 3</intersection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-178.5,27.5,-178</points>
<connection>
<GID>554</GID>
<name>OUT_0</name></connection>
<intersection>-178 2</intersection></vsegment></shape></wire>
<wire>
<ID>660 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-154.5,-39,-154.5</points>
<connection>
<GID>504</GID>
<name>IN_1</name></connection>
<connection>
<GID>510</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>325 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-101.5,-29,-89</points>
<intersection>-101.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,-89,-29,-89</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29,-101.5,-26.5,-101.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>335 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-103.5,-30,-99</points>
<intersection>-103.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-103.5,-26.5,-103.5</points>
<connection>
<GID>233</GID>
<name>IN_3</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-99,-30,-99</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>346 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-119,-29,-107.5</points>
<intersection>-119 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-107.5,-26.5,-107.5</points>
<connection>
<GID>233</GID>
<name>IN_4</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-119,-29,-119</points>
<connection>
<GID>288</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>343 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-114,-29.5,-106.5</points>
<intersection>-114 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-106.5,-26.5,-106.5</points>
<connection>
<GID>233</GID>
<name>IN_5</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-114,-29.5,-114</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>338 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-104.5,-30,-104</points>
<intersection>-104.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-104.5,-26.5,-104.5</points>
<connection>
<GID>233</GID>
<name>IN_7</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-104,-30,-104</points>
<connection>
<GID>272</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>331 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-104,-18.5,-104</points>
<connection>
<GID>233</GID>
<name>OUT</name></connection>
<connection>
<GID>258</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>633 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-149.5,16,-149.5</points>
<connection>
<GID>475</GID>
<name>IN_1</name></connection>
<connection>
<GID>482</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>328 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-88,-39,-88</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>327 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-90,-39,-90</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<connection>
<GID>248</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>497 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-110,126,-110</points>
<connection>
<GID>394</GID>
<name>IN_1</name></connection>
<connection>
<GID>401</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>704 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-187.5,16,-187.5</points>
<connection>
<GID>570</GID>
<name>IN_0</name></connection>
<connection>
<GID>571</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>856 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-223.5,-30,-223</points>
<intersection>-223.5 1</intersection>
<intersection>-223 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-223.5,-26.5,-223.5</points>
<connection>
<GID>704</GID>
<name>IN_7</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-223,-30,-223</points>
<connection>
<GID>715</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>711 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-189.5,16,-189.5</points>
<connection>
<GID>570</GID>
<name>IN_1</name></connection>
<connection>
<GID>575</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>703 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-188.5,25,-185</points>
<intersection>-188.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-185,28.5,-185</points>
<connection>
<GID>556</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-188.5,25,-188.5</points>
<connection>
<GID>570</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>330 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-91,-53,-91</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-55,-105,-55,-91</points>
<intersection>-105 6</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-55,-105,-53,-105</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment></shape></wire>
<wire>
<ID>693 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-170.5,2,-170.5</points>
<connection>
<GID>558</GID>
<name>IN_1</name></connection>
<connection>
<GID>561</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>0,-184.5,0,-170.5</points>
<intersection>-184.5 6</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>0,-184.5,2,-184.5</points>
<connection>
<GID>568</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment></shape></wire>
<wire>
<ID>637 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-141,-29,-128.5</points>
<intersection>-141 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,-128.5,-29,-128.5</points>
<connection>
<GID>489</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29,-141,-26.5,-141</points>
<connection>
<GID>488</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>332 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-93,-39,-93</points>
<connection>
<GID>262</GID>
<name>IN_0</name></connection>
<connection>
<GID>260</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>699 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-177.5,16,-177.5</points>
<connection>
<GID>565</GID>
<name>IN_0</name></connection>
<connection>
<GID>566</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>692 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-168.5,2,-168.5</points>
<connection>
<GID>558</GID>
<name>IN_0</name></connection>
<connection>
<GID>560</GID>
<name>IN_0</name></connection>
<intersection>1 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1,-179.5,1,-168.5</points>
<intersection>-179.5 8</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>1,-179.5,16,-179.5</points>
<connection>
<GID>565</GID>
<name>IN_1</name></connection>
<intersection>1 7</intersection></hsegment></shape></wire>
<wire>
<ID>698 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-183,25,-178.5</points>
<intersection>-183 1</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-183,28.5,-183</points>
<connection>
<GID>556</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-178.5,25,-178.5</points>
<connection>
<GID>565</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>702 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-182.5,16,-182.5</points>
<connection>
<GID>569</GID>
<name>IN_0</name></connection>
<connection>
<GID>567</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>336 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-98,-39,-98</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<connection>
<GID>268</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>706 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-192.5,16,-192.5</points>
<connection>
<GID>573</GID>
<name>IN_0</name></connection>
<connection>
<GID>572</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>340 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-103,-39,-103</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<connection>
<GID>276</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>339 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-105,-39,-105</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<connection>
<GID>274</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>342 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-108,-39,-108</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>415 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-110,-39,-110</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<connection>
<GID>318</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>344 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-113,-39,-113</points>
<connection>
<GID>282</GID>
<name>IN_0</name></connection>
<connection>
<GID>284</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>416 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-115,-39,-115</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<connection>
<GID>320</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>772 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145.5,-223,146.5,-223</points>
<connection>
<GID>626</GID>
<name>OUT</name></connection>
<connection>
<GID>625</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>617 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-132.5,16,-132.5</points>
<connection>
<GID>468</GID>
<name>IN_0</name></connection>
<connection>
<GID>467</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>440 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-100.5,28.5,-98.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-98.5,28.5,-98.5</points>
<intersection>27.5 3</intersection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-99,27.5,-98.5</points>
<connection>
<GID>324</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>769 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-207,126,-207</points>
<connection>
<GID>629</GID>
<name>IN_0</name></connection>
<connection>
<GID>627</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>601 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-153.5,80.5,-146</points>
<intersection>-153.5 2</intersection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-146,83.5,-146</points>
<connection>
<GID>434</GID>
<name>IN_5</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-153.5,80.5,-153.5</points>
<connection>
<GID>450</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>424 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-104,36.5,-104</points>
<connection>
<GID>326</GID>
<name>OUT</name></connection>
<connection>
<GID>325</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>419 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-101.5,26,-89</points>
<intersection>-101.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-89,26,-89</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-101.5,28.5,-101.5</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>427 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-102.5,25.5,-94</points>
<intersection>-102.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-102.5,28.5,-102.5</points>
<connection>
<GID>326</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-94,25.5,-94</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>605 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-159.5,71,-159.5</points>
<connection>
<GID>453</GID>
<name>IN_1</name></connection>
<connection>
<GID>454</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>428 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-103.5,25,-99</points>
<intersection>-103.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-103.5,28.5,-103.5</points>
<connection>
<GID>326</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-99,25,-99</points>
<connection>
<GID>335</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>438 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-119,26,-107.5</points>
<intersection>-119 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-107.5,28.5,-107.5</points>
<connection>
<GID>326</GID>
<name>IN_4</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-119,26,-119</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>435 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-114,25.5,-106.5</points>
<intersection>-114 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-106.5,28.5,-106.5</points>
<connection>
<GID>326</GID>
<name>IN_5</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-114,25.5,-114</points>
<connection>
<GID>342</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>640 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-128.5,-53,-128.5</points>
<connection>
<GID>490</GID>
<name>IN_0</name></connection>
<connection>
<GID>492</GID>
<name>IN_0</name></connection>
<intersection>-54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-54,-139.5,-54,-128.5</points>
<intersection>-139.5 8</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-54,-139.5,-39,-139.5</points>
<connection>
<GID>497</GID>
<name>IN_1</name></connection>
<intersection>-54 7</intersection></hsegment></shape></wire>
<wire>
<ID>433 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-109,25,-105.5</points>
<intersection>-109 2</intersection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-105.5,28.5,-105.5</points>
<connection>
<GID>326</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-109,25,-109</points>
<connection>
<GID>340</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>430 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-104.5,25,-104</points>
<intersection>-104.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-104.5,28.5,-104.5</points>
<connection>
<GID>326</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-104,25,-104</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>756 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-187.5,126,-187.5</points>
<connection>
<GID>613</GID>
<name>IN_0</name></connection>
<connection>
<GID>614</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>421 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-88,16,-88</points>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<connection>
<GID>327</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>420 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-90,16,-90</points>
<connection>
<GID>328</GID>
<name>OUT</name></connection>
<connection>
<GID>327</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>422 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-89,2,-89</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<intersection>1 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1,-100,1,-89</points>
<intersection>-100 8</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>1,-100,16,-100</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>1 7</intersection></hsegment></shape></wire>
<wire>
<ID>423 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-91,2,-91</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>0,-105,0,-91</points>
<intersection>-105 6</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>0,-105,2,-105</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment></shape></wire>
<wire>
<ID>773 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-212,126,-212</points>
<connection>
<GID>633</GID>
<name>IN_0</name></connection>
<connection>
<GID>632</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>653 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-153.5,-29.5,-146</points>
<intersection>-153.5 2</intersection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-146,-26.5,-146</points>
<connection>
<GID>488</GID>
<name>IN_5</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-153.5,-29.5,-153.5</points>
<connection>
<GID>504</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>476 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145.5,-104,146.5,-104</points>
<connection>
<GID>380</GID>
<name>OUT</name></connection>
<connection>
<GID>379</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>806 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-222,71,-222</points>
<connection>
<GID>664</GID>
<name>IN_0</name></connection>
<connection>
<GID>666</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>467 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-110,71,-110</points>
<connection>
<GID>367</GID>
<name>IN_1</name></connection>
<connection>
<GID>374</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>805 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-224,71,-224</points>
<connection>
<GID>664</GID>
<name>IN_1</name></connection>
<connection>
<GID>665</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>643 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-132.5,-39,-132.5</points>
<connection>
<GID>495</GID>
<name>IN_0</name></connection>
<connection>
<GID>494</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>804 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-223.5,80,-223</points>
<intersection>-223.5 1</intersection>
<intersection>-223 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-223.5,83.5,-223.5</points>
<connection>
<GID>653</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-223,80,-223</points>
<connection>
<GID>664</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>425 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-93,16,-93</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<connection>
<GID>332</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>426 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-95,16,-95</points>
<connection>
<GID>332</GID>
<name>IN_1</name></connection>
<connection>
<GID>334</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>747 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-172.5,126,-172.5</points>
<connection>
<GID>605</GID>
<name>IN_0</name></connection>
<connection>
<GID>606</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>780 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-222,126,-222</points>
<connection>
<GID>637</GID>
<name>IN_0</name></connection>
<connection>
<GID>639</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>657 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-159.5,-39,-159.5</points>
<connection>
<GID>507</GID>
<name>IN_1</name></connection>
<connection>
<GID>508</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>480 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-103.5,135,-99</points>
<intersection>-103.5 1</intersection>
<intersection>-99 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-103.5,138.5,-103.5</points>
<connection>
<GID>380</GID>
<name>IN_3</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-99,135,-99</points>
<connection>
<GID>389</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>810 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-232,71,-232</points>
<connection>
<GID>668</GID>
<name>IN_0</name></connection>
<connection>
<GID>669</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>809 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-233,80.5,-225.5</points>
<intersection>-233 2</intersection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-225.5,83.5,-225.5</points>
<connection>
<GID>653</GID>
<name>IN_5</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-233,80.5,-233</points>
<connection>
<GID>668</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>764 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-194.5,126,-194.5</points>
<connection>
<GID>615</GID>
<name>IN_1</name></connection>
<connection>
<GID>621</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>429 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-98,16,-98</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<connection>
<GID>335</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>432 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-103,16,-103</points>
<connection>
<GID>339</GID>
<name>IN_0</name></connection>
<connection>
<GID>337</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>431 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-105,16,-105</points>
<connection>
<GID>338</GID>
<name>OUT_0</name></connection>
<connection>
<GID>337</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>434 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-108,16,-108</points>
<connection>
<GID>341</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>648 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-144,-30,-143.5</points>
<intersection>-144 1</intersection>
<intersection>-143.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-144,-26.5,-144</points>
<connection>
<GID>488</GID>
<name>IN_7</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-143.5,-30,-143.5</points>
<connection>
<GID>499</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>441 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-110,16,-110</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<connection>
<GID>347</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>613 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-127.5,16,-127.5</points>
<connection>
<GID>464</GID>
<name>IN_0</name></connection>
<connection>
<GID>462</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>436 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-113,16,-113</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<connection>
<GID>342</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>442 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-115,16,-115</points>
<connection>
<GID>342</GID>
<name>IN_1</name></connection>
<connection>
<GID>348</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>483 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-105,126,-105</points>
<connection>
<GID>392</GID>
<name>OUT_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>821 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-207,16,-207</points>
<connection>
<GID>680</GID>
<name>IN_0</name></connection>
<connection>
<GID>682</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>659 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-149.5,-39,-149.5</points>
<connection>
<GID>502</GID>
<name>IN_1</name></connection>
<connection>
<GID>509</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>820 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-209,16,-209</points>
<connection>
<GID>680</GID>
<name>IN_1</name></connection>
<connection>
<GID>681</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>819 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-220.5,26,-208</points>
<intersection>-220.5 2</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-208,26,-208</points>
<connection>
<GID>680</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-220.5,28.5,-220.5</points>
<connection>
<GID>679</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>852 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-214,-39,-214</points>
<connection>
<GID>710</GID>
<name>IN_1</name></connection>
<connection>
<GID>712</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>853 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-221.5,-29.5,-213</points>
<intersection>-221.5 1</intersection>
<intersection>-213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-221.5,-26.5,-221.5</points>
<connection>
<GID>704</GID>
<name>IN_2</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-213,-29.5,-213</points>
<connection>
<GID>710</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>503 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-127.5,126,-127.5</points>
<connection>
<GID>410</GID>
<name>IN_0</name></connection>
<connection>
<GID>408</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>825 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-212,16,-212</points>
<connection>
<GID>684</GID>
<name>IN_0</name></connection>
<connection>
<GID>685</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>827 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-221.5,25.5,-213</points>
<intersection>-221.5 1</intersection>
<intersection>-213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-221.5,28.5,-221.5</points>
<connection>
<GID>679</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-213,25.5,-213</points>
<connection>
<GID>684</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>631 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-159.5,16,-159.5</points>
<connection>
<GID>480</GID>
<name>IN_1</name></connection>
<connection>
<GID>481</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>466 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-100.5,83.5,-98.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<intersection>-98.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-98.5,83.5,-98.5</points>
<intersection>82.5 3</intersection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-99,82.5,-98.5</points>
<connection>
<GID>351</GID>
<name>OUT_0</name></connection>
<intersection>-98.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>453 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-102.5,80.5,-94</points>
<intersection>-102.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-102.5,83.5,-102.5</points>
<connection>
<GID>353</GID>
<name>IN_2</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-94,80.5,-94</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>461 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-114,80.5,-106.5</points>
<intersection>-114 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-106.5,83.5,-106.5</points>
<connection>
<GID>353</GID>
<name>IN_5</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-114,80.5,-114</points>
<connection>
<GID>369</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>797 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-210,57,-210</points>
<connection>
<GID>655</GID>
<name>IN_1</name></connection>
<connection>
<GID>658</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>55,-224,55,-210</points>
<intersection>-224 6</intersection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>55,-224,57,-224</points>
<connection>
<GID>665</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment></shape></wire>
<wire>
<ID>459 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-109,80,-105.5</points>
<intersection>-109 2</intersection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-105.5,83.5,-105.5</points>
<connection>
<GID>353</GID>
<name>IN_6</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-109,80,-109</points>
<connection>
<GID>367</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>491 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-114,135.5,-106.5</points>
<intersection>-114 2</intersection>
<intersection>-106.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-106.5,138.5,-106.5</points>
<connection>
<GID>380</GID>
<name>IN_5</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-114,135.5,-114</points>
<connection>
<GID>396</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>829 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-217,16,-217</points>
<connection>
<GID>688</GID>
<name>IN_0</name></connection>
<connection>
<GID>687</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>449 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-91,57,-91</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>55,-105,55,-91</points>
<intersection>-105 6</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>55,-105,57,-105</points>
<connection>
<GID>365</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment></shape></wire>
<wire>
<ID>860 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-227,-39,-227</points>
<connection>
<GID>718</GID>
<name>IN_0</name></connection>
<connection>
<GID>719</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>859 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-228,-30,-224.5</points>
<intersection>-228 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-224.5,-26.5,-224.5</points>
<connection>
<GID>704</GID>
<name>IN_6</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-228,-30,-228</points>
<connection>
<GID>718</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>834 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-227,16,-227</points>
<connection>
<GID>692</GID>
<name>IN_0</name></connection>
<connection>
<GID>693</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>841 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-229,16,-229</points>
<connection>
<GID>692</GID>
<name>IN_1</name></connection>
<connection>
<GID>699</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>833 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-228,25,-224.5</points>
<intersection>-228 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-224.5,28.5,-224.5</points>
<connection>
<GID>679</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-228,25,-228</points>
<connection>
<GID>692</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>757 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-193.5,135.5,-186</points>
<intersection>-193.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-186,138.5,-186</points>
<connection>
<GID>599</GID>
<name>IN_5</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-193.5,135.5,-193.5</points>
<connection>
<GID>615</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>782 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-227,126,-227</points>
<connection>
<GID>640</GID>
<name>IN_0</name></connection>
<connection>
<GID>641</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>452 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-95,71,-95</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<connection>
<GID>361</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>848 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-208,-53,-208</points>
<connection>
<GID>706</GID>
<name>IN_0</name></connection>
<connection>
<GID>708</GID>
<name>IN_0</name></connection>
<intersection>-54 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-54,-219,-54,-208</points>
<intersection>-219 8</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-54,-219,-39,-219</points>
<connection>
<GID>713</GID>
<name>IN_1</name></connection>
<intersection>-54 7</intersection></hsegment></shape></wire>
<wire>
<ID>849 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-56,-210,-53,-210</points>
<connection>
<GID>706</GID>
<name>IN_1</name></connection>
<connection>
<GID>709</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-55,-224,-55,-210</points>
<intersection>-224 6</intersection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-55,-224,-53,-224</points>
<connection>
<GID>716</GID>
<name>IN_0</name></connection>
<intersection>-55 5</intersection></hsegment></shape></wire>
<wire>
<ID>846 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-209,-39,-209</points>
<connection>
<GID>706</GID>
<name>OUT</name></connection>
<connection>
<GID>705</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>868 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-234,-39,-234</points>
<connection>
<GID>720</GID>
<name>IN_1</name></connection>
<connection>
<GID>726</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>842 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-234,16,-234</points>
<connection>
<GID>694</GID>
<name>IN_1</name></connection>
<connection>
<GID>700</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>790 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-234,126,-234</points>
<connection>
<GID>642</GID>
<name>IN_1</name></connection>
<connection>
<GID>648</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>460 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-108,71,-108</points>
<connection>
<GID>368</GID>
<name>IN_0</name></connection>
<connection>
<GID>367</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>855 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-217,-39,-217</points>
<connection>
<GID>714</GID>
<name>IN_0</name></connection>
<connection>
<GID>713</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>686 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-194.5,-39,-194.5</points>
<connection>
<GID>545</GID>
<name>IN_1</name></connection>
<connection>
<GID>551</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>611 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-141,26,-128.5</points>
<intersection>-141 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-128.5,26,-128.5</points>
<connection>
<GID>462</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-141,28.5,-141</points>
<connection>
<GID>461</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>462 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-113,71,-113</points>
<connection>
<GID>370</GID>
<name>IN_0</name></connection>
<connection>
<GID>369</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>645 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-142,-29.5,-133.5</points>
<intersection>-142 1</intersection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-142,-26.5,-142</points>
<connection>
<GID>488</GID>
<name>IN_2</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-133.5,-29.5,-133.5</points>
<connection>
<GID>494</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>798 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-223,91.5,-223</points>
<connection>
<GID>653</GID>
<name>OUT</name></connection>
<connection>
<GID>652</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>468 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-115,71,-115</points>
<connection>
<GID>369</GID>
<name>IN_1</name></connection>
<connection>
<GID>375</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>505 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-130.5,112,-130.5</points>
<connection>
<GID>409</GID>
<name>IN_1</name></connection>
<connection>
<GID>412</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>110,-144.5,110,-130.5</points>
<intersection>-144.5 6</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>110,-144.5,112,-144.5</points>
<connection>
<GID>419</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment></shape></wire>
<wire>
<ID>712 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-194.5,16,-194.5</points>
<connection>
<GID>572</GID>
<name>IN_1</name></connection>
<connection>
<GID>576</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>873 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-188,82.5,-187</points>
<connection>
<GID>734</GID>
<name>OUT_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-187,83.5,-187</points>
<connection>
<GID>579</GID>
<name>IN_4</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>718 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-168.5,57,-168.5</points>
<connection>
<GID>580</GID>
<name>IN_0</name></connection>
<connection>
<GID>581</GID>
<name>IN_0</name></connection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>56,-179.5,56,-168.5</points>
<intersection>-179.5 8</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>56,-179.5,71,-179.5</points>
<connection>
<GID>524</GID>
<name>IN_1</name></connection>
<intersection>56 7</intersection></hsegment></shape></wire>
<wire>
<ID>719 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-170.5,57,-170.5</points>
<connection>
<GID>580</GID>
<name>IN_1</name></connection>
<connection>
<GID>582</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>55,-184.5,55,-170.5</points>
<intersection>-184.5 6</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>55,-184.5,57,-184.5</points>
<connection>
<GID>586</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment></shape></wire>
<wire>
<ID>509 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-142,135.5,-133.5</points>
<intersection>-142 1</intersection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-142,138.5,-142</points>
<connection>
<GID>407</GID>
<name>IN_2</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-133.5,135.5,-133.5</points>
<connection>
<GID>413</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>716 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-169.5,71,-169.5</points>
<connection>
<GID>580</GID>
<name>OUT</name></connection>
<connection>
<GID>514</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>722 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-174.5,71,-174.5</points>
<connection>
<GID>583</GID>
<name>IN_1</name></connection>
<connection>
<GID>584</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>877 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,-227.5,82.5,-226.5</points>
<connection>
<GID>742</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-226.5,83.5,-226.5</points>
<connection>
<GID>653</GID>
<name>IN_4</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>793 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-220.5,81,-208</points>
<intersection>-220.5 2</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-208,81,-208</points>
<connection>
<GID>654</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-220.5,83.5,-220.5</points>
<connection>
<GID>653</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>471 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-101.5,136,-89</points>
<intersection>-101.5 2</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-89,136,-89</points>
<connection>
<GID>381</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>136,-101.5,138.5,-101.5</points>
<connection>
<GID>380</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>801 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-221.5,80.5,-213</points>
<intersection>-221.5 1</intersection>
<intersection>-213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-221.5,83.5,-221.5</points>
<connection>
<GID>653</GID>
<name>IN_2</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-213,80.5,-213</points>
<connection>
<GID>659</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>479 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-102.5,135.5,-94</points>
<intersection>-102.5 1</intersection>
<intersection>-94 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-102.5,138.5,-102.5</points>
<connection>
<GID>380</GID>
<name>IN_2</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-94,135.5,-94</points>
<connection>
<GID>386</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>494 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-119,136,-107.5</points>
<intersection>-119 2</intersection>
<intersection>-107.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>136,-107.5,138.5,-107.5</points>
<connection>
<GID>380</GID>
<name>IN_4</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-119,136,-119</points>
<connection>
<GID>399</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>485 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-109,135,-105.5</points>
<intersection>-109 2</intersection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-105.5,138.5,-105.5</points>
<connection>
<GID>380</GID>
<name>IN_6</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-109,135,-109</points>
<connection>
<GID>394</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>482 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-104.5,135,-104</points>
<intersection>-104.5 1</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-104.5,138.5,-104.5</points>
<connection>
<GID>380</GID>
<name>IN_7</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-104,135,-104</points>
<connection>
<GID>391</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>691 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-167.5,16,-167.5</points>
<connection>
<GID>557</GID>
<name>IN_0</name></connection>
<connection>
<GID>559</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>690 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-169.5,16,-169.5</points>
<connection>
<GID>557</GID>
<name>IN_1</name></connection>
<connection>
<GID>558</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>689 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-181,26,-168.5</points>
<intersection>-181 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>22,-168.5,26,-168.5</points>
<connection>
<GID>557</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26,-181,28.5,-181</points>
<connection>
<GID>556</GID>
<name>IN_1</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>473 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-88,126,-88</points>
<connection>
<GID>383</GID>
<name>IN_0</name></connection>
<connection>
<GID>381</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>649 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-144.5,-39,-144.5</points>
<connection>
<GID>500</GID>
<name>OUT_0</name></connection>
<connection>
<GID>499</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>802 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-222.5,80,-218</points>
<intersection>-222.5 1</intersection>
<intersection>-218 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-222.5,83.5,-222.5</points>
<connection>
<GID>653</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-218,80,-218</points>
<connection>
<GID>662</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>472 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-90,126,-90</points>
<connection>
<GID>382</GID>
<name>OUT</name></connection>
<connection>
<GID>381</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>730 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-187.5,71,-187.5</points>
<connection>
<GID>588</GID>
<name>IN_0</name></connection>
<connection>
<GID>587</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>639 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-127.5,-39,-127.5</points>
<connection>
<GID>491</GID>
<name>IN_0</name></connection>
<connection>
<GID>489</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>474 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-89,112,-89</points>
<connection>
<GID>382</GID>
<name>IN_0</name></connection>
<connection>
<GID>384</GID>
<name>IN_0</name></connection>
<intersection>111 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-100,111,-89</points>
<intersection>-100 8</intersection>
<intersection>-89 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>111,-100,126,-100</points>
<connection>
<GID>389</GID>
<name>IN_1</name></connection>
<intersection>111 7</intersection></hsegment></shape></wire>
<wire>
<ID>475 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-91,112,-91</points>
<connection>
<GID>382</GID>
<name>IN_1</name></connection>
<connection>
<GID>385</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>110,-105,110,-91</points>
<intersection>-105 6</intersection>
<intersection>-91 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>110,-105,112,-105</points>
<connection>
<GID>392</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment></shape></wire>
<wire>
<ID>832 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-222,16,-222</points>
<connection>
<GID>689</GID>
<name>IN_0</name></connection>
<connection>
<GID>691</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>831 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-224,16,-224</points>
<connection>
<GID>689</GID>
<name>IN_1</name></connection>
<connection>
<GID>690</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>862 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-232,-39,-232</points>
<connection>
<GID>720</GID>
<name>IN_0</name></connection>
<connection>
<GID>721</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>861 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29.5,-233,-29.5,-225.5</points>
<intersection>-233 2</intersection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29.5,-225.5,-26.5,-225.5</points>
<connection>
<GID>704</GID>
<name>IN_5</name></connection>
<intersection>-29.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-233,-29.5,-233</points>
<connection>
<GID>720</GID>
<name>OUT</name></connection>
<intersection>-29.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>477 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-93,126,-93</points>
<connection>
<GID>387</GID>
<name>IN_0</name></connection>
<connection>
<GID>386</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>627 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-153.5,25.5,-146</points>
<intersection>-153.5 2</intersection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-146,28.5,-146</points>
<connection>
<GID>461</GID>
<name>IN_5</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-153.5,25.5,-153.5</points>
<connection>
<GID>477</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>478 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-95,126,-95</points>
<connection>
<GID>386</GID>
<name>IN_1</name></connection>
<connection>
<GID>388</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>481 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-98,126,-98</points>
<connection>
<GID>390</GID>
<name>IN_0</name></connection>
<connection>
<GID>389</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>814 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-219.5,83.5,-217.5</points>
<connection>
<GID>653</GID>
<name>IN_0</name></connection>
<intersection>-217.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-217.5,83.5,-217.5</points>
<intersection>82.5 3</intersection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-218,82.5,-217.5</points>
<connection>
<GID>651</GID>
<name>OUT_0</name></connection>
<intersection>-217.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>484 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-103,126,-103</points>
<connection>
<GID>393</GID>
<name>IN_0</name></connection>
<connection>
<GID>391</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>527 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-152.5,126,-152.5</points>
<connection>
<GID>424</GID>
<name>IN_0</name></connection>
<connection>
<GID>423</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>490 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-108,126,-108</points>
<connection>
<GID>395</GID>
<name>IN_0</name></connection>
<connection>
<GID>394</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>822 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-208,2,-208</points>
<connection>
<GID>681</GID>
<name>IN_0</name></connection>
<connection>
<GID>516</GID>
<name>IN_0</name></connection>
<intersection>1 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>1,-219,1,-208</points>
<intersection>-219 8</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>1,-219,16,-219</points>
<connection>
<GID>687</GID>
<name>IN_1</name></connection>
<intersection>1 7</intersection></hsegment></shape></wire>
<wire>
<ID>669 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-172.5,-39,-172.5</points>
<connection>
<GID>535</GID>
<name>IN_0</name></connection>
<connection>
<GID>536</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>492 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-113,126,-113</points>
<connection>
<GID>397</GID>
<name>IN_0</name></connection>
<connection>
<GID>396</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>498 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-115,126,-115</points>
<connection>
<GID>396</GID>
<name>IN_1</name></connection>
<connection>
<GID>402</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>493 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>125,-118,126,-118</points>
<connection>
<GID>398</GID>
<name>IN_0</name></connection>
<connection>
<GID>399</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>495 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-120,126,-120</points>
<connection>
<GID>399</GID>
<name>IN_1</name></connection>
<connection>
<GID>400</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>721 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-172.5,71,-172.5</points>
<connection>
<GID>527</GID>
<name>IN_0</name></connection>
<connection>
<GID>583</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>874 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-188,137.5,-187</points>
<connection>
<GID>736</GID>
<name>OUT_0</name></connection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-187,138.5,-187</points>
<connection>
<GID>599</GID>
<name>IN_4</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>701 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-184.5,16,-184.5</points>
<connection>
<GID>567</GID>
<name>IN_1</name></connection>
<connection>
<GID>568</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>700 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-184,25,-183.5</points>
<intersection>-184 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-184,28.5,-184</points>
<connection>
<GID>556</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-183.5,25,-183.5</points>
<connection>
<GID>567</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>510 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-143,135,-138.5</points>
<intersection>-143 1</intersection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-143,138.5,-143</points>
<connection>
<GID>407</GID>
<name>IN_3</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-138.5,135,-138.5</points>
<connection>
<GID>416</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>531 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-140,138.5,-138</points>
<connection>
<GID>407</GID>
<name>IN_0</name></connection>
<intersection>-138 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-138,138.5,-138</points>
<intersection>137.5 3</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>137.5,-138.5,137.5,-138</points>
<connection>
<GID>405</GID>
<name>OUT_0</name></connection>
<intersection>-138 2</intersection></vsegment></shape></wire>
<wire>
<ID>715 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-181,81,-168.5</points>
<intersection>-181 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-168.5,81,-168.5</points>
<connection>
<GID>514</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-181,83.5,-181</points>
<connection>
<GID>579</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>876 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,-227.5,27.5,-226.5</points>
<connection>
<GID>740</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,-226.5,28.5,-226.5</points>
<connection>
<GID>679</GID>
<name>IN_4</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>506 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145.5,-143.5,146.5,-143.5</points>
<connection>
<GID>407</GID>
<name>OUT</name></connection>
<connection>
<GID>406</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>694 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-183.5,36.5,-183.5</points>
<connection>
<GID>556</GID>
<name>OUT</name></connection>
<connection>
<GID>555</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>501 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-141,136,-128.5</points>
<intersection>-141 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-128.5,136,-128.5</points>
<connection>
<GID>408</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>136,-141,138.5,-141</points>
<connection>
<GID>407</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>526 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-153.5,135.5,-146</points>
<intersection>-153.5 2</intersection>
<intersection>-146 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-146,138.5,-146</points>
<connection>
<GID>407</GID>
<name>IN_5</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-153.5,135.5,-153.5</points>
<connection>
<GID>423</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>524 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-148.5,135,-145</points>
<intersection>-148.5 2</intersection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-145,138.5,-145</points>
<connection>
<GID>407</GID>
<name>IN_6</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-148.5,135,-148.5</points>
<connection>
<GID>421</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>523 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-142.5,126,-142.5</points>
<connection>
<GID>420</GID>
<name>IN_0</name></connection>
<connection>
<GID>418</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>502 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-129.5,126,-129.5</points>
<connection>
<GID>409</GID>
<name>OUT</name></connection>
<connection>
<GID>408</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>878 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-227.5,137.5,-226.5</points>
<connection>
<GID>744</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-226.5,138.5,-226.5</points>
<connection>
<GID>626</GID>
<name>IN_4</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>725 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-177.5,71,-177.5</points>
<connection>
<GID>585</GID>
<name>IN_0</name></connection>
<connection>
<GID>524</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>504 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-128.5,112,-128.5</points>
<connection>
<GID>409</GID>
<name>IN_0</name></connection>
<connection>
<GID>411</GID>
<name>IN_0</name></connection>
<intersection>111 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-139.5,111,-128.5</points>
<intersection>-139.5 8</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>111,-139.5,126,-139.5</points>
<connection>
<GID>416</GID>
<name>IN_1</name></connection>
<intersection>111 7</intersection></hsegment></shape></wire>
<wire>
<ID>732 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-192.5,71,-192.5</points>
<connection>
<GID>589</GID>
<name>IN_0</name></connection>
<connection>
<GID>590</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>731 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-193.5,80.5,-186</points>
<intersection>-193.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-186,83.5,-186</points>
<connection>
<GID>579</GID>
<name>IN_5</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-193.5,80.5,-193.5</points>
<connection>
<GID>589</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>507 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-132.5,126,-132.5</points>
<connection>
<GID>414</GID>
<name>IN_0</name></connection>
<connection>
<GID>413</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>695 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-172.5,16,-172.5</points>
<connection>
<GID>563</GID>
<name>IN_0</name></connection>
<connection>
<GID>562</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>511 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-137.5,126,-137.5</points>
<connection>
<GID>417</GID>
<name>IN_0</name></connection>
<connection>
<GID>416</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>737 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-189.5,71,-189.5</points>
<connection>
<GID>587</GID>
<name>IN_1</name></connection>
<connection>
<GID>593</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>522 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116,-144.5,126,-144.5</points>
<connection>
<GID>419</GID>
<name>OUT_0</name></connection>
<connection>
<GID>418</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>762 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-180,138.5,-178</points>
<connection>
<GID>599</GID>
<name>IN_0</name></connection>
<intersection>-178 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-178,138.5,-178</points>
<intersection>137.5 3</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>137.5,-178.5,137.5,-178</points>
<connection>
<GID>597</GID>
<name>OUT_0</name></connection>
<intersection>-178 2</intersection></vsegment></shape></wire>
<wire>
<ID>532 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-149.5,126,-149.5</points>
<connection>
<GID>421</GID>
<name>IN_1</name></connection>
<connection>
<GID>428</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>533 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-154.5,126,-154.5</points>
<connection>
<GID>423</GID>
<name>IN_1</name></connection>
<connection>
<GID>429</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>744 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-168.5,112,-168.5</points>
<connection>
<GID>601</GID>
<name>IN_0</name></connection>
<connection>
<GID>603</GID>
<name>IN_0</name></connection>
<intersection>111 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-179.5,111,-168.5</points>
<intersection>-179.5 8</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>111,-179.5,126,-179.5</points>
<connection>
<GID>608</GID>
<name>IN_1</name></connection>
<intersection>111 7</intersection></hsegment></shape></wire>
<wire>
<ID>770 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-208,112,-208</points>
<connection>
<GID>628</GID>
<name>IN_0</name></connection>
<connection>
<GID>630</GID>
<name>IN_0</name></connection>
<intersection>111 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>111,-219,111,-208</points>
<intersection>-219 8</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>111,-219,126,-219</points>
<connection>
<GID>635</GID>
<name>IN_1</name></connection>
<intersection>111 7</intersection></hsegment></shape></wire>
<wire>
<ID>745 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-170.5,112,-170.5</points>
<connection>
<GID>601</GID>
<name>IN_1</name></connection>
<connection>
<GID>604</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>110,-184.5,110,-170.5</points>
<intersection>-184.5 6</intersection>
<intersection>-170.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>110,-184.5,112,-184.5</points>
<connection>
<GID>611</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment></shape></wire>
<wire>
<ID>742 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-169.5,126,-169.5</points>
<connection>
<GID>601</GID>
<name>OUT</name></connection>
<connection>
<GID>600</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>528 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-157.5,126,-157.5</points>
<connection>
<GID>426</GID>
<name>IN_0</name></connection>
<connection>
<GID>425</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>530 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-159.5,126,-159.5</points>
<connection>
<GID>426</GID>
<name>IN_1</name></connection>
<connection>
<GID>427</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>748 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-174.5,126,-174.5</points>
<connection>
<GID>605</GID>
<name>IN_1</name></connection>
<connection>
<GID>607</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>774 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-214,126,-214</points>
<connection>
<GID>632</GID>
<name>IN_1</name></connection>
<connection>
<GID>634</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>749 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-182,135.5,-173.5</points>
<intersection>-182 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-182,138.5,-182</points>
<connection>
<GID>599</GID>
<name>IN_2</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-173.5,135.5,-173.5</points>
<connection>
<GID>605</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>606 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-140,83.5,-138</points>
<connection>
<GID>434</GID>
<name>IN_0</name></connection>
<intersection>-138 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-138,83.5,-138</points>
<intersection>82.5 3</intersection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-138.5,82.5,-138</points>
<connection>
<GID>432</GID>
<name>OUT_0</name></connection>
<intersection>-138 2</intersection></vsegment></shape></wire>
<wire>
<ID>768 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-209,126,-209</points>
<connection>
<GID>627</GID>
<name>IN_1</name></connection>
<connection>
<GID>628</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>751 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-177.5,126,-177.5</points>
<connection>
<GID>609</GID>
<name>IN_0</name></connection>
<connection>
<GID>608</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>541 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-143.5,91.5,-143.5</points>
<connection>
<GID>434</GID>
<name>OUT</name></connection>
<connection>
<GID>433</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>781 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-228,135,-224.5</points>
<intersection>-228 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-224.5,138.5,-224.5</points>
<connection>
<GID>626</GID>
<name>IN_6</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-228,135,-228</points>
<connection>
<GID>640</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>536 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-141,81,-128.5</points>
<intersection>-141 2</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-128.5,81,-128.5</points>
<connection>
<GID>435</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-141,83.5,-141</points>
<connection>
<GID>434</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>586 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-142,80.5,-133.5</points>
<intersection>-142 1</intersection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-142,83.5,-142</points>
<connection>
<GID>434</GID>
<name>IN_2</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-133.5,80.5,-133.5</points>
<connection>
<GID>440</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>587 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-143,80,-138.5</points>
<intersection>-143 1</intersection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-143,83.5,-143</points>
<connection>
<GID>434</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-138.5,80,-138.5</points>
<connection>
<GID>443</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>599 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-148.5,80,-145</points>
<intersection>-148.5 2</intersection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-145,83.5,-145</points>
<connection>
<GID>434</GID>
<name>IN_6</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-148.5,80,-148.5</points>
<connection>
<GID>448</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>589 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-144,80,-143.5</points>
<intersection>-144 1</intersection>
<intersection>-143.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-144,83.5,-144</points>
<connection>
<GID>434</GID>
<name>IN_7</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-143.5,80,-143.5</points>
<connection>
<GID>445</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>537 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,-129.5,71,-129.5</points>
<connection>
<GID>436</GID>
<name>OUT</name></connection>
<connection>
<GID>435</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>539 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-128.5,57,-128.5</points>
<connection>
<GID>436</GID>
<name>IN_0</name></connection>
<connection>
<GID>438</GID>
<name>IN_0</name></connection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>56,-139.5,56,-128.5</points>
<intersection>-139.5 8</intersection>
<intersection>-128.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>56,-139.5,71,-139.5</points>
<connection>
<GID>443</GID>
<name>IN_1</name></connection>
<intersection>56 7</intersection></hsegment></shape></wire>
<wire>
<ID>540 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-130.5,57,-130.5</points>
<connection>
<GID>436</GID>
<name>IN_1</name></connection>
<connection>
<GID>439</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>55,-144.5,55,-130.5</points>
<intersection>-144.5 6</intersection>
<intersection>-130.5 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>55,-144.5,57,-144.5</points>
<connection>
<GID>446</GID>
<name>IN_0</name></connection>
<intersection>55 5</intersection></hsegment></shape></wire>
<wire>
<ID>796 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-208,57,-208</points>
<connection>
<GID>655</GID>
<name>IN_0</name></connection>
<connection>
<GID>657</GID>
<name>IN_0</name></connection>
<intersection>56 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>56,-219,56,-208</points>
<intersection>-219 8</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>56,-219,71,-219</points>
<connection>
<GID>662</GID>
<name>IN_1</name></connection>
<intersection>56 7</intersection></hsegment></shape></wire>
<wire>
<ID>763 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-189.5,126,-189.5</points>
<connection>
<GID>613</GID>
<name>IN_1</name></connection>
<connection>
<GID>620</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>788 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138.5,-219.5,138.5,-217.5</points>
<connection>
<GID>626</GID>
<name>IN_0</name></connection>
<intersection>-217.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-217.5,138.5,-217.5</points>
<intersection>137.5 3</intersection>
<intersection>138.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>137.5,-218,137.5,-217.5</points>
<connection>
<GID>624</GID>
<name>OUT_0</name></connection>
<intersection>-217.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>755 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-188.5,135,-185</points>
<intersection>-188.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-185,138.5,-185</points>
<connection>
<GID>599</GID>
<name>IN_6</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-188.5,135,-188.5</points>
<connection>
<GID>613</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>579 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-132.5,71,-132.5</points>
<connection>
<GID>441</GID>
<name>IN_0</name></connection>
<connection>
<GID>440</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>585 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-134.5,71,-134.5</points>
<connection>
<GID>440</GID>
<name>IN_1</name></connection>
<connection>
<GID>442</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>588 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-137.5,71,-137.5</points>
<connection>
<GID>444</GID>
<name>IN_0</name></connection>
<connection>
<GID>443</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>598 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-142.5,71,-142.5</points>
<connection>
<GID>447</GID>
<name>IN_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>590 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,-144.5,71,-144.5</points>
<connection>
<GID>446</GID>
<name>OUT_0</name></connection>
<connection>
<GID>445</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>607 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-149.5,71,-149.5</points>
<connection>
<GID>448</GID>
<name>IN_1</name></connection>
<connection>
<GID>455</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>602 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-152.5,71,-152.5</points>
<connection>
<GID>451</GID>
<name>IN_0</name></connection>
<connection>
<GID>450</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>616 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-143.5,36.5,-143.5</points>
<connection>
<GID>461</GID>
<name>OUT</name></connection>
<connection>
<GID>460</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>619 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-142,25.5,-133.5</points>
<intersection>-142 1</intersection>
<intersection>-133.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-142,28.5,-142</points>
<connection>
<GID>461</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-133.5,25.5,-133.5</points>
<connection>
<GID>467</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>620 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-143,25,-138.5</points>
<intersection>-143 1</intersection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-143,28.5,-143</points>
<connection>
<GID>461</GID>
<name>IN_3</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-138.5,25,-138.5</points>
<connection>
<GID>470</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>630 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-158.5,26,-147</points>
<intersection>-158.5 2</intersection>
<intersection>-147 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-147,28.5,-147</points>
<connection>
<GID>461</GID>
<name>IN_4</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-158.5,26,-158.5</points>
<connection>
<GID>480</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>625 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-148.5,25,-145</points>
<intersection>-148.5 2</intersection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-145,28.5,-145</points>
<connection>
<GID>461</GID>
<name>IN_6</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-148.5,25,-148.5</points>
<connection>
<GID>475</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>622 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-144,25,-143.5</points>
<intersection>-144 1</intersection>
<intersection>-143.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25,-144,28.5,-144</points>
<connection>
<GID>461</GID>
<name>IN_7</name></connection>
<intersection>25 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-143.5,25,-143.5</points>
<connection>
<GID>472</GID>
<name>OUT</name></connection>
<intersection>25 0</intersection></hsegment></shape></wire>
<wire>
<ID>612 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>8,-129.5,16,-129.5</points>
<connection>
<GID>463</GID>
<name>OUT</name></connection>
<connection>
<GID>462</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>771 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>109,-210,112,-210</points>
<connection>
<GID>628</GID>
<name>IN_1</name></connection>
<connection>
<GID>631</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>110,-224,110,-210</points>
<intersection>-224 6</intersection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>110,-224,112,-224</points>
<connection>
<GID>638</GID>
<name>IN_0</name></connection>
<intersection>110 5</intersection></hsegment></shape></wire>
<wire>
<ID>618 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-134.5,16,-134.5</points>
<connection>
<GID>467</GID>
<name>IN_1</name></connection>
<connection>
<GID>469</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>621 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-137.5,16,-137.5</points>
<connection>
<GID>471</GID>
<name>IN_0</name></connection>
<connection>
<GID>470</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>624 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-142.5,16,-142.5</points>
<connection>
<GID>474</GID>
<name>IN_0</name></connection>
<connection>
<GID>472</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>626 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-147.5,16,-147.5</points>
<connection>
<GID>476</GID>
<name>IN_0</name></connection>
<connection>
<GID>475</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>807 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-228,80,-224.5</points>
<intersection>-228 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-224.5,83.5,-224.5</points>
<connection>
<GID>653</GID>
<name>IN_6</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-228,80,-228</points>
<connection>
<GID>667</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>634 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-154.5,16,-154.5</points>
<connection>
<GID>477</GID>
<name>IN_1</name></connection>
<connection>
<GID>483</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>784 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-232,126,-232</points>
<connection>
<GID>642</GID>
<name>IN_0</name></connection>
<connection>
<GID>643</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>767 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-220.5,136,-208</points>
<intersection>-220.5 2</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-208,136,-208</points>
<connection>
<GID>627</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>136,-220.5,138.5,-220.5</points>
<connection>
<GID>626</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>629 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-157.5,16,-157.5</points>
<connection>
<GID>479</GID>
<name>IN_0</name></connection>
<connection>
<GID>480</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>655 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-157.5,-39,-157.5</points>
<connection>
<GID>506</GID>
<name>IN_0</name></connection>
<connection>
<GID>507</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>800 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-214,71,-214</points>
<connection>
<GID>659</GID>
<name>IN_1</name></connection>
<connection>
<GID>661</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>658 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-140,-26.5,-138</points>
<connection>
<GID>488</GID>
<name>IN_0</name></connection>
<intersection>-138 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-138,-26.5,-138</points>
<intersection>-27.5 3</intersection>
<intersection>-26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-138.5,-27.5,-138</points>
<connection>
<GID>486</GID>
<name>OUT_0</name></connection>
<intersection>-138 2</intersection></vsegment></shape></wire>
<wire>
<ID>776 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-222.5,135,-218</points>
<intersection>-222.5 1</intersection>
<intersection>-218 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-222.5,138.5,-222.5</points>
<connection>
<GID>626</GID>
<name>IN_3</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-218,135,-218</points>
<connection>
<GID>635</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>646 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-143,-30,-138.5</points>
<intersection>-143 1</intersection>
<intersection>-138.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-143,-26.5,-143</points>
<connection>
<GID>488</GID>
<name>IN_3</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-138.5,-30,-138.5</points>
<connection>
<GID>497</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>656 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-158.5,-29,-147</points>
<intersection>-158.5 2</intersection>
<intersection>-147 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-29,-147,-26.5,-147</points>
<connection>
<GID>488</GID>
<name>IN_4</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-158.5,-29,-158.5</points>
<connection>
<GID>507</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>651 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-148.5,-30,-145</points>
<intersection>-148.5 2</intersection>
<intersection>-145 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-145,-26.5,-145</points>
<connection>
<GID>488</GID>
<name>IN_6</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-148.5,-30,-148.5</points>
<connection>
<GID>502</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>638 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-47,-129.5,-39,-129.5</points>
<connection>
<GID>490</GID>
<name>OUT</name></connection>
<connection>
<GID>489</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>815 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-229,71,-229</points>
<connection>
<GID>667</GID>
<name>IN_1</name></connection>
<connection>
<GID>673</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>647 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-137.5,-39,-137.5</points>
<connection>
<GID>498</GID>
<name>IN_0</name></connection>
<connection>
<GID>497</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>866 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,-219.5,-26.5,-217.5</points>
<connection>
<GID>704</GID>
<name>IN_0</name></connection>
<intersection>-217.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,-217.5,-26.5,-217.5</points>
<intersection>-27.5 3</intersection>
<intersection>-26.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-27.5,-218,-27.5,-217.5</points>
<connection>
<GID>702</GID>
<name>OUT_0</name></connection>
<intersection>-217.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>845 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-29,-220.5,-29,-208</points>
<intersection>-220.5 2</intersection>
<intersection>-208 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,-208,-29,-208</points>
<connection>
<GID>705</GID>
<name>OUT</name></connection>
<intersection>-29 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-29,-220.5,-26.5,-220.5</points>
<connection>
<GID>704</GID>
<name>IN_1</name></connection>
<intersection>-29 0</intersection></hsegment></shape></wire>
<wire>
<ID>854 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,-222.5,-30,-218</points>
<intersection>-222.5 1</intersection>
<intersection>-218 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-30,-222.5,-26.5,-222.5</points>
<connection>
<GID>704</GID>
<name>IN_3</name></connection>
<intersection>-30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-218,-30,-218</points>
<connection>
<GID>713</GID>
<name>OUT</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>875 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-27.5,-227.5,-27.5,-226.5</points>
<connection>
<GID>738</GID>
<name>OUT_0</name></connection>
<intersection>-226.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,-226.5,-26.5,-226.5</points>
<connection>
<GID>704</GID>
<name>IN_4</name></connection>
<intersection>-27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>850 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19.5,-223,-18.5,-223</points>
<connection>
<GID>704</GID>
<name>OUT</name></connection>
<connection>
<GID>703</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>840 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-219.5,28.5,-217.5</points>
<connection>
<GID>679</GID>
<name>IN_0</name></connection>
<intersection>-217.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>27.5,-217.5,28.5,-217.5</points>
<intersection>27.5 3</intersection>
<intersection>28.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>27.5,-218,27.5,-217.5</points>
<connection>
<GID>677</GID>
<name>OUT_0</name></connection>
<intersection>-217.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>720 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-183.5,91.5,-183.5</points>
<connection>
<GID>579</GID>
<name>OUT</name></connection>
<connection>
<GID>523</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>823 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-1,-210,2,-210</points>
<connection>
<GID>681</GID>
<name>IN_1</name></connection>
<connection>
<GID>683</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>0,-224,0,-210</points>
<intersection>-224 6</intersection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>0,-224,2,-224</points>
<connection>
<GID>690</GID>
<name>IN_0</name></connection>
<intersection>0 5</intersection></hsegment></shape></wire>
<wire>
<ID>678 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-187.5,-39,-187.5</points>
<connection>
<GID>543</GID>
<name>IN_0</name></connection>
<connection>
<GID>544</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>857 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-49,-224,-39,-224</points>
<connection>
<GID>716</GID>
<name>OUT_0</name></connection>
<connection>
<GID>715</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>717 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-167.5,71,-167.5</points>
<connection>
<GID>514</GID>
<name>IN_0</name></connection>
<connection>
<GID>520</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>724 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-183,80,-178.5</points>
<intersection>-183 1</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-183,83.5,-183</points>
<connection>
<GID>579</GID>
<name>IN_3</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-178.5,80,-178.5</points>
<connection>
<GID>524</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>697 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-182,25.5,-173.5</points>
<intersection>-182 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-182,28.5,-182</points>
<connection>
<GID>556</GID>
<name>IN_2</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-173.5,25.5,-173.5</points>
<connection>
<GID>562</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>858 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-222,-39,-222</points>
<connection>
<GID>715</GID>
<name>IN_0</name></connection>
<connection>
<GID>717</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>705 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-193.5,25.5,-186</points>
<intersection>-193.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-186,28.5,-186</points>
<connection>
<GID>556</GID>
<name>IN_5</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-193.5,25.5,-193.5</points>
<connection>
<GID>572</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>696 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-174.5,16,-174.5</points>
<connection>
<GID>562</GID>
<name>IN_1</name></connection>
<connection>
<GID>564</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>736 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-180,83.5,-178</points>
<connection>
<GID>579</GID>
<name>IN_0</name></connection>
<intersection>-178 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-178,83.5,-178</points>
<intersection>82.5 3</intersection>
<intersection>83.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-178.5,82.5,-178</points>
<connection>
<GID>578</GID>
<name>OUT_0</name></connection>
<intersection>-178 2</intersection></vsegment></shape></wire>
<wire>
<ID>723 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80.5,-182,80.5,-173.5</points>
<intersection>-182 1</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80.5,-182,83.5,-182</points>
<connection>
<GID>579</GID>
<name>IN_2</name></connection>
<intersection>80.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-173.5,80.5,-173.5</points>
<connection>
<GID>583</GID>
<name>OUT</name></connection>
<intersection>80.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>729 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-188.5,80,-185</points>
<intersection>-188.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>80,-185,83.5,-185</points>
<connection>
<GID>579</GID>
<name>IN_6</name></connection>
<intersection>80 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>77,-188.5,80,-188.5</points>
<connection>
<GID>587</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>741 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>136,-181,136,-168.5</points>
<intersection>-181 2</intersection>
<intersection>-168.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>132,-168.5,136,-168.5</points>
<connection>
<GID>600</GID>
<name>OUT</name></connection>
<intersection>136 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>136,-181,138.5,-181</points>
<connection>
<GID>599</GID>
<name>IN_1</name></connection>
<intersection>136 0</intersection></hsegment></shape></wire>
<wire>
<ID>752 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135,-184,135,-183.5</points>
<intersection>-184 1</intersection>
<intersection>-183.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135,-184,138.5,-184</points>
<connection>
<GID>599</GID>
<name>IN_7</name></connection>
<intersection>135 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-183.5,135,-183.5</points>
<connection>
<GID>610</GID>
<name>OUT</name></connection>
<intersection>135 0</intersection></hsegment></shape></wire>
<wire>
<ID>743 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-167.5,126,-167.5</points>
<connection>
<GID>600</GID>
<name>IN_0</name></connection>
<connection>
<GID>602</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>754 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>125,-182.5,126,-182.5</points>
<connection>
<GID>610</GID>
<name>IN_0</name></connection>
<connection>
<GID>612</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>775 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-221.5,135.5,-213</points>
<intersection>-221.5 1</intersection>
<intersection>-213 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-221.5,138.5,-221.5</points>
<connection>
<GID>626</GID>
<name>IN_2</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-213,135.5,-213</points>
<connection>
<GID>632</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>783 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-233,135.5,-225.5</points>
<intersection>-233 2</intersection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-225.5,138.5,-225.5</points>
<connection>
<GID>626</GID>
<name>IN_5</name></connection>
<intersection>135.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132,-233,135.5,-233</points>
<connection>
<GID>642</GID>
<name>OUT</name></connection>
<intersection>135.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>795 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-207,71,-207</points>
<connection>
<GID>654</GID>
<name>IN_0</name></connection>
<connection>
<GID>656</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>803 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-217,71,-217</points>
<connection>
<GID>662</GID>
<name>IN_0</name></connection>
<connection>
<GID>663</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>835 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25.5,-233,25.5,-225.5</points>
<intersection>-233 2</intersection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>25.5,-225.5,28.5,-225.5</points>
<connection>
<GID>679</GID>
<name>IN_5</name></connection>
<intersection>25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22,-233,25.5,-233</points>
<connection>
<GID>694</GID>
<name>OUT</name></connection>
<intersection>25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>836 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-232,16,-232</points>
<connection>
<GID>694</GID>
<name>IN_0</name></connection>
<connection>
<GID>695</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>847 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-207,-39,-207</points>
<connection>
<GID>705</GID>
<name>IN_0</name></connection>
<connection>
<GID>707</GID>
<name>IN_0</name></connection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-154.475,141.592,152.95,-13.6752</PageViewport>
<gate>
<ID>754</ID>
<type>DA_FROM</type>
<position>127,17</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR10</lparam></gate>
<gate>
<ID>279</ID>
<type>DA_FROM</type>
<position>-73,85</position>
<input>
<ID>IN_0</ID>337 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>168</ID>
<type>DE_TO</type>
<position>-10.5,52</position>
<input>
<ID>IN_0</ID>636 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>232</ID>
<type>DE_TO</type>
<position>-15,24</position>
<input>
<ID>IN_0</ID>408 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T8</lparam></gate>
<gate>
<ID>921</ID>
<type>DA_FROM</type>
<position>72.5,69.5</position>
<input>
<ID>IN_0</ID>1039 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC=0</lparam></gate>
<gate>
<ID>160</ID>
<type>DE_TO</type>
<position>-16,51</position>
<input>
<ID>IN_0</ID>609 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>849</ID>
<type>DA_FROM</type>
<position>-118,84.5</position>
<input>
<ID>IN_0</ID>950 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo12</lparam></gate>
<gate>
<ID>779</ID>
<type>DA_FROM</type>
<position>18,50</position>
<input>
<ID>IN_0</ID>923 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>246</ID>
<type>DE_TO</type>
<position>-10.5,54</position>
<input>
<ID>IN_0</ID>683 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>748</ID>
<type>DE_TO</type>
<position>-61,117</position>
<input>
<ID>IN_0</ID>959 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AND</lparam></gate>
<gate>
<ID>917</ID>
<type>DA_FROM</type>
<position>72.5,78.5</position>
<input>
<ID>IN_0</ID>1043 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR3</lparam></gate>
<gate>
<ID>228</ID>
<type>DE_TO</type>
<position>-15,22</position>
<input>
<ID>IN_0</ID>361 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>259</ID>
<type>DE_TO</type>
<position>-61,95</position>
<input>
<ID>IN_0</ID>322 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIR</lparam></gate>
<gate>
<ID>750</ID>
<type>DE_TO</type>
<position>-61,111.5</position>
<input>
<ID>IN_0</ID>964 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ADD</lparam></gate>
<gate>
<ID>323</ID>
<type>DA_FROM</type>
<position>-78,62</position>
<input>
<ID>IN_0</ID>1132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR15</lparam></gate>
<gate>
<ID>49</ID>
<type>AA_AND2</type>
<position>-131,50.5</position>
<input>
<ID>IN_0</ID>80 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>78 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>751</ID>
<type>DA_FROM</type>
<position>65.5,125.5</position>
<input>
<ID>IN_0</ID>896 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>768</ID>
<type>DE_TO</type>
<position>37,66</position>
<input>
<ID>IN_0</ID>1103 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mem_W</lparam></gate>
<gate>
<ID>58</ID>
<type>DA_FROM</type>
<position>10,10</position>
<input>
<ID>IN_0</ID>16 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>752</ID>
<type>DE_TO</type>
<position>-61,106</position>
<input>
<ID>IN_0</ID>999 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID LDA</lparam></gate>
<gate>
<ID>175</ID>
<type>DE_TO</type>
<position>-8.5,19</position>
<input>
<ID>IN_0</ID>355 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>756</ID>
<type>AA_LABEL</type>
<position>134.5,23.5</position>
<gparam>LABEL_TEXT Output Register Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>10,2</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /I</lparam></gate>
<gate>
<ID>925</ID>
<type>AE_OR4</type>
<position>16,33.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<input>
<ID>IN_1</ID>1097 </input>
<input>
<ID>IN_2</ID>1098 </input>
<input>
<ID>IN_3</ID>1099 </input>
<output>
<ID>OUT</ID>1095 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>236</ID>
<type>DE_TO</type>
<position>-8.5,27</position>
<input>
<ID>IN_0</ID>353 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T11</lparam></gate>
<gate>
<ID>1040</ID>
<type>DA_FROM</type>
<position>-78.5,12.5</position>
<input>
<ID>IN_0</ID>904 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>172</ID>
<type>DE_TO</type>
<position>-15,16</position>
<input>
<ID>IN_0</ID>411 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>759</ID>
<type>DA_FROM</type>
<position>-78.5,17.5</position>
<input>
<ID>IN_0</ID>1143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>776</ID>
<type>BE_NOR2</type>
<position>-104,108</position>
<input>
<ID>IN_0</ID>910 </input>
<input>
<ID>IN_1</ID>911 </input>
<output>
<ID>OUT</ID>934 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>DA_FROM</type>
<position>10,12</position>
<input>
<ID>IN_0</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>994</ID>
<type>DA_FROM</type>
<position>-78.5,40.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_REGISTER4</type>
<position>-31,17</position>
<output>
<ID>OUT_0</ID>77 </output>
<output>
<ID>OUT_1</ID>204 </output>
<output>
<ID>OUT_2</ID>191 </output>
<output>
<ID>OUT_3</ID>203 </output>
<input>
<ID>clear</ID>242 </input>
<input>
<ID>clock</ID>205 </input>
<input>
<ID>count_enable</ID>319 </input>
<gparam>VALUE_BOX -0.8,-0.8,0.8,1.8</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>MAX_COUNT 15</lparam>
<lparam>SYNC_CLEAR true</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>815</ID>
<type>AE_OR3</type>
<position>31,44</position>
<input>
<ID>IN_0</ID>942 </input>
<input>
<ID>IN_1</ID>1100 </input>
<input>
<ID>IN_2</ID>941 </input>
<output>
<ID>OUT</ID>939 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>138</ID>
<type>BI_DECODER_4x16</type>
<position>-23,23.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>204 </input>
<input>
<ID>IN_2</ID>191 </input>
<input>
<ID>IN_3</ID>203 </input>
<output>
<ID>OUT_0</ID>411 </output>
<output>
<ID>OUT_1</ID>359 </output>
<output>
<ID>OUT_10</ID>407 </output>
<output>
<ID>OUT_11</ID>353 </output>
<output>
<ID>OUT_12</ID>410 </output>
<output>
<ID>OUT_13</ID>354 </output>
<output>
<ID>OUT_14</ID>412 </output>
<output>
<ID>OUT_15</ID>356 </output>
<output>
<ID>OUT_2</ID>406 </output>
<output>
<ID>OUT_3</ID>355 </output>
<output>
<ID>OUT_4</ID>409 </output>
<output>
<ID>OUT_5</ID>357 </output>
<output>
<ID>OUT_6</ID>361 </output>
<output>
<ID>OUT_7</ID>358 </output>
<output>
<ID>OUT_8</ID>408 </output>
<output>
<ID>OUT_9</ID>360 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>803</ID>
<type>DE_TO</type>
<position>-98,108</position>
<input>
<ID>IN_0</ID>934 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR=0</lparam></gate>
<gate>
<ID>142</ID>
<type>DA_FROM</type>
<position>-35.5,11.5</position>
<input>
<ID>IN_0</ID>205 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>833</ID>
<type>DA_FROM</type>
<position>-28,118</position>
<input>
<ID>IN_0</ID>1078 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>144</ID>
<type>DA_FROM</type>
<position>-35.5,9.5</position>
<input>
<ID>IN_0</ID>242 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SCclr</lparam></gate>
<gate>
<ID>823</ID>
<type>DA_FROM</type>
<position>-118,94.5</position>
<input>
<ID>IN_0</ID>967 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo2</lparam></gate>
<gate>
<ID>146</ID>
<type>DA_FROM</type>
<position>-35,24</position>
<input>
<ID>IN_0</ID>319 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s</lparam></gate>
<gate>
<ID>148</ID>
<type>AA_AND2</type>
<position>133,18</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>837</ID>
<type>DA_FROM</type>
<position>-127.5,89.5</position>
<input>
<ID>IN_0</ID>1006 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo7</lparam></gate>
<gate>
<ID>1003</ID>
<type>DA_FROM</type>
<position>-89,39.5</position>
<input>
<ID>IN_0</ID>1175 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR8</lparam></gate>
<gate>
<ID>317</ID>
<type>DA_FROM</type>
<position>-69,57.5</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>152</ID>
<type>DA_FROM</type>
<position>118,102</position>
<input>
<ID>IN_0</ID>898 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>841</ID>
<type>AA_AND2</type>
<position>-67,111.5</position>
<input>
<ID>IN_0</ID>962 </input>
<input>
<ID>IN_1</ID>963 </input>
<output>
<ID>OUT</ID>964 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1026</ID>
<type>AA_AND4</type>
<position>-72.5,37.5</position>
<input>
<ID>IN_0</ID>1173 </input>
<input>
<ID>IN_1</ID>1174 </input>
<input>
<ID>IN_2</ID>1193 </input>
<input>
<ID>IN_3</ID>1194 </input>
<output>
<ID>OUT</ID>1201 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>158</ID>
<type>BE_JKFF_LOW</type>
<position>-63,57.5</position>
<input>
<ID>J</ID>1130 </input>
<input>
<ID>K</ID>1131 </input>
<output>
<ID>Q</ID>886 </output>
<input>
<ID>clock</ID>23 </input>
<output>
<ID>nQ</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>819</ID>
<type>AA_AND2</type>
<position>80,19</position>
<input>
<ID>IN_0</ID>1180 </input>
<input>
<ID>IN_1</ID>1179 </input>
<output>
<ID>OUT</ID>948 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>DE_TO</type>
<position>-15,28</position>
<input>
<ID>IN_0</ID>410 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T12</lparam></gate>
<gate>
<ID>1041</ID>
<type>DA_FROM</type>
<position>-89,11.5</position>
<input>
<ID>IN_0</ID>938 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR8</lparam></gate>
<gate>
<ID>1020</ID>
<type>AE_OR2</type>
<position>-65,29.5</position>
<input>
<ID>IN_0</ID>1155 </input>
<input>
<ID>IN_1</ID>1201 </input>
<output>
<ID>OUT</ID>1153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>DE_TO</type>
<position>-8.5,17</position>
<input>
<ID>IN_0</ID>359 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>46</ID>
<type>BE_DECODER_3x8</type>
<position>-23,50.5</position>
<input>
<ID>IN_0</ID>534 </input>
<input>
<ID>IN_1</ID>500 </input>
<input>
<ID>IN_2</ID>499 </input>
<output>
<ID>OUT_0</ID>610 </output>
<output>
<ID>OUT_1</ID>661 </output>
<output>
<ID>OUT_2</ID>635 </output>
<output>
<ID>OUT_3</ID>682 </output>
<output>
<ID>OUT_4</ID>609 </output>
<output>
<ID>OUT_5</ID>636 </output>
<output>
<ID>OUT_6</ID>535 </output>
<output>
<ID>OUT_7</ID>683 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>771</ID>
<type>DA_FROM</type>
<position>18,43</position>
<input>
<ID>IN_0</ID>1101 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>238</ID>
<type>DE_TO</type>
<position>-8.5,29</position>
<input>
<ID>IN_0</ID>354 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T13</lparam></gate>
<gate>
<ID>1042</ID>
<type>DA_FROM</type>
<position>-89,9.5</position>
<input>
<ID>IN_0</ID>1010 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>174</ID>
<type>DE_TO</type>
<position>-15,18</position>
<input>
<ID>IN_0</ID>406 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>283</ID>
<type>DA_FROM</type>
<position>-73,83</position>
<input>
<ID>IN_0</ID>349 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR11</lparam></gate>
<gate>
<ID>646</ID>
<type>DE_TO</type>
<position>85,114</position>
<input>
<ID>IN_0</ID>1035 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_CLR</lparam></gate>
<gate>
<ID>877</ID>
<type>DA_FROM</type>
<position>-89,1.5</position>
<input>
<ID>IN_0</ID>1159 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR6</lparam></gate>
<gate>
<ID>1056</ID>
<type>AA_AND2</type>
<position>80,10</position>
<input>
<ID>IN_0</ID>1187 </input>
<input>
<ID>IN_1</ID>1184 </input>
<output>
<ID>OUT</ID>1183 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>DE_TO</type>
<position>-15,20</position>
<input>
<ID>IN_0</ID>409 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>988</ID>
<type>DA_FROM</type>
<position>-86,58.5</position>
<input>
<ID>IN_0</ID>1135 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>294</ID>
<type>DE_TO</type>
<position>-109.5,-0.5</position>
<input>
<ID>IN_0</ID>351 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>141</ID>
<type>DA_FROM</type>
<position>-29.5,48</position>
<input>
<ID>IN_0</ID>500 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR13</lparam></gate>
<gate>
<ID>205</ID>
<type>DE_TO</type>
<position>-8.5,21</position>
<input>
<ID>IN_0</ID>357 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>891</ID>
<type>DA_FROM</type>
<position>125.5,54</position>
<input>
<ID>IN_0</ID>1089 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>230</ID>
<type>DE_TO</type>
<position>-8.5,23</position>
<input>
<ID>IN_0</ID>358 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T7</lparam></gate>
<gate>
<ID>234</ID>
<type>DE_TO</type>
<position>-8.5,25</position>
<input>
<ID>IN_0</ID>360 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T9</lparam></gate>
<gate>
<ID>783</ID>
<type>AE_SMALL_INVERTER</type>
<position>-15.5,56.5</position>
<input>
<ID>IN_0</ID>683 </input>
<output>
<ID>OUT_0</ID>914 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>170</ID>
<type>DE_TO</type>
<position>-16,53</position>
<input>
<ID>IN_0</ID>535 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>235</ID>
<type>DE_TO</type>
<position>-15,26</position>
<input>
<ID>IN_0</ID>407 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T10</lparam></gate>
<gate>
<ID>791</ID>
<type>DA_FROM</type>
<position>-126,106.5</position>
<input>
<ID>IN_0</ID>929 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR9</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_TO</type>
<position>-15,30</position>
<input>
<ID>IN_0</ID>412 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T14</lparam></gate>
<gate>
<ID>933</ID>
<type>AA_AND2</type>
<position>65,57.5</position>
<input>
<ID>IN_0</ID>1054 </input>
<input>
<ID>IN_1</ID>1053 </input>
<output>
<ID>OUT</ID>1052 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>574</ID>
<type>DA_FROM</type>
<position>18,105</position>
<input>
<ID>IN_0</ID>791 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>244</ID>
<type>DE_TO</type>
<position>-8.5,31</position>
<input>
<ID>IN_0</ID>356 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T15</lparam></gate>
<gate>
<ID>83</ID>
<type>DA_FROM</type>
<position>-29.5,46</position>
<input>
<ID>IN_0</ID>534 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR12</lparam></gate>
<gate>
<ID>1031</ID>
<type>DA_FROM</type>
<position>-78.5,48.5</position>
<input>
<ID>IN_0</ID>1163 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>147</ID>
<type>DE_TO</type>
<position>-16,47</position>
<input>
<ID>IN_0</ID>610 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>308</ID>
<type>GA_LED</type>
<position>-112.5,62</position>
<input>
<ID>N_in2</ID>733 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>143</ID>
<type>DA_FROM</type>
<position>-29.5,50</position>
<input>
<ID>IN_0</ID>499 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR14</lparam></gate>
<gate>
<ID>996</ID>
<type>AE_SMALL_INVERTER</type>
<position>-14.5,11</position>
<input>
<ID>IN_0</ID>359 </input>
<output>
<ID>OUT_0</ID>1138 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>149</ID>
<type>DE_TO</type>
<position>-10.5,48</position>
<input>
<ID>IN_0</ID>661 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>302</ID>
<type>BE_JKFF_LOW</type>
<position>-116.5,57.5</position>
<input>
<ID>J</ID>1127 </input>
<input>
<ID>K</ID>75 </input>
<output>
<ID>Q</ID>733 </output>
<input>
<ID>clock</ID>470 </input>
<output>
<ID>nQ</ID>469 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>-16,49</position>
<input>
<ID>IN_0</ID>635 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>296</ID>
<type>DA_FROM</type>
<position>-64,26</position>
<input>
<ID>IN_0</ID>443 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>1000</ID>
<type>DE_TO</type>
<position>-11,9</position>
<input>
<ID>IN_0</ID>1139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /T2</lparam></gate>
<gate>
<ID>153</ID>
<type>DE_TO</type>
<position>-10.5,50</position>
<input>
<ID>IN_0</ID>682 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>306</ID>
<type>DE_TO</type>
<position>-109.5,59.5</position>
<input>
<ID>IN_0</ID>733 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IEN</lparam></gate>
<gate>
<ID>321</ID>
<type>DE_TO</type>
<position>-56,59.5</position>
<input>
<ID>IN_0</ID>886 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>592</ID>
<type>DE_TO</type>
<position>37,109</position>
<input>
<ID>IN_0</ID>954 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_CLR</lparam></gate>
<gate>
<ID>257</ID>
<type>DA_FROM</type>
<position>-73,99.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR9</lparam></gate>
<gate>
<ID>762</ID>
<type>DE_TO</type>
<position>137.5,34</position>
<input>
<ID>IN_0</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_CLR</lparam></gate>
<gate>
<ID>287</ID>
<type>DA_FROM</type>
<position>-122.5,1.5</position>
<input>
<ID>IN_0</ID>352 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>553</ID>
<type>DE_TO</type>
<position>37,100</position>
<input>
<ID>IN_0</ID>882 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_INC</lparam></gate>
<gate>
<ID>376</ID>
<type>AA_AND2</type>
<position>24,126</position>
<input>
<ID>IN_0</ID>734 </input>
<input>
<ID>IN_1</ID>740 </input>
<output>
<ID>OUT</ID>739 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>577</ID>
<type>DE_TO</type>
<position>37,124</position>
<input>
<ID>IN_0</ID>735 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_LD</lparam></gate>
<gate>
<ID>596</ID>
<type>DE_TO</type>
<position>37,89.5</position>
<input>
<ID>IN_0</ID>883 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AR_bus</lparam></gate>
<gate>
<ID>261</ID>
<type>DA_FROM</type>
<position>-73,96</position>
<input>
<ID>IN_0</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>981</ID>
<type>AE_SMALL_INVERTER</type>
<position>-89,4.5</position>
<input>
<ID>IN_0</ID>1161 </input>
<output>
<ID>OUT_0</ID>1160 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>622</ID>
<type>DE_TO</type>
<position>107.5,82</position>
<input>
<ID>IN_0</ID>1008 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_INC</lparam></gate>
<gate>
<ID>644</ID>
<type>DE_TO</type>
<position>84.5,126.5</position>
<input>
<ID>IN_0</ID>900 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_LD</lparam></gate>
<gate>
<ID>650</ID>
<type>DE_TO</type>
<position>84.5,44.5</position>
<input>
<ID>IN_0</ID>1067 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID PC_bus</lparam></gate>
<gate>
<ID>303</ID>
<type>DE_TO</type>
<position>-109.5,42</position>
<input>
<ID>IN_0</ID>687 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /FGI</lparam></gate>
<gate>
<ID>698</ID>
<type>DE_TO</type>
<position>137.5,110.5</position>
<input>
<ID>IN_0</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_INC</lparam></gate>
<gate>
<ID>701</ID>
<type>DE_TO</type>
<position>137.5,128</position>
<input>
<ID>IN_0</ID>930 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_LD</lparam></gate>
<gate>
<ID>1060</ID>
<type>DA_FROM</type>
<position>62,10</position>
<input>
<ID>IN_0</ID>1185 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>722</ID>
<type>DE_TO</type>
<position>137.5,99</position>
<input>
<ID>IN_0</ID>1009 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_bus</lparam></gate>
<gate>
<ID>872</ID>
<type>DA_FROM</type>
<position>-73,107</position>
<input>
<ID>IN_0</ID>997 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>727</ID>
<type>DE_TO</type>
<position>-10,85</position>
<input>
<ID>IN_0</ID>1081 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_CLR</lparam></gate>
<gate>
<ID>728</ID>
<type>DE_TO</type>
<position>-10,91</position>
<input>
<ID>IN_0</ID>1064 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_INC</lparam></gate>
<gate>
<ID>1059</ID>
<type>DA_FROM</type>
<position>62,8</position>
<input>
<ID>IN_0</ID>1186 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>882</ID>
<type>DA_FROM</type>
<position>-22,90</position>
<input>
<ID>IN_0</ID>1079 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR5</lparam></gate>
<gate>
<ID>729</ID>
<type>DE_TO</type>
<position>-9,113</position>
<input>
<ID>IN_0</ID>1017 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_LD</lparam></gate>
<gate>
<ID>892</ID>
<type>AA_AND2</type>
<position>131.5,53</position>
<input>
<ID>IN_0</ID>1089 </input>
<input>
<ID>IN_1</ID>1090 </input>
<output>
<ID>OUT</ID>1091 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>731</ID>
<type>DE_TO</type>
<position>-10,77</position>
<input>
<ID>IN_0</ID>1087 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC_bus</lparam></gate>
<gate>
<ID>735</ID>
<type>DE_TO</type>
<position>137.5,74.5</position>
<input>
<ID>IN_0</ID>1013 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR_LD</lparam></gate>
<gate>
<ID>880</ID>
<type>DE_OR8</type>
<position>100.5,82</position>
<input>
<ID>IN_0</ID>1026 </input>
<input>
<ID>IN_1</ID>1025 </input>
<input>
<ID>IN_2</ID>1024 </input>
<input>
<ID>IN_3</ID>1023 </input>
<input>
<ID>IN_4</ID>1019 </input>
<input>
<ID>IN_5</ID>1020 </input>
<input>
<ID>IN_6</ID>1021 </input>
<input>
<ID>IN_7</ID>1022 </input>
<output>
<ID>OUT</ID>1008 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1067</ID>
<type>DA_FROM</type>
<position>74,4.5</position>
<input>
<ID>IN_0</ID>1189 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>890</ID>
<type>FF_GND</type>
<position>134,39.5</position>
<output>
<ID>OUT_0</ID>1088 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>737</ID>
<type>DE_TO</type>
<position>137.5,69</position>
<input>
<ID>IN_0</ID>1016 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR_bus</lparam></gate>
<gate>
<ID>745</ID>
<type>DA_FROM</type>
<position>-35,107.5</position>
<input>
<ID>IN_0</ID>24 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR6</lparam></gate>
<gate>
<ID>770</ID>
<type>DE_OR8</type>
<position>-112,112</position>
<input>
<ID>IN_0</ID>912 </input>
<input>
<ID>IN_1</ID>924 </input>
<input>
<ID>IN_2</ID>916 </input>
<input>
<ID>IN_3</ID>926 </input>
<input>
<ID>IN_4</ID>921 </input>
<input>
<ID>IN_5</ID>915 </input>
<input>
<ID>IN_6</ID>927 </input>
<input>
<ID>IN_7</ID>913 </input>
<output>
<ID>OUT</ID>910 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>1075</ID>
<type>AE_OR2</type>
<position>-16,85</position>
<input>
<ID>IN_0</ID>1129 </input>
<input>
<ID>IN_1</ID>1084 </input>
<output>
<ID>OUT</ID>1081 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>761</ID>
<type>AA_AND2</type>
<position>-22,100.5</position>
<input>
<ID>IN_0</ID>1072 </input>
<input>
<ID>IN_1</ID>1071 </input>
<output>
<ID>OUT</ID>1070 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>786</ID>
<type>DA_FROM</type>
<position>-118,111.5</position>
<input>
<ID>IN_0</ID>913 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR4</lparam></gate>
<gate>
<ID>763</ID>
<type>DE_TO</type>
<position>137.5,41.5</position>
<input>
<ID>IN_0</ID>1088 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_INC</lparam></gate>
<gate>
<ID>796</ID>
<type>DA_FROM</type>
<position>-118,103.5</position>
<input>
<ID>IN_0</ID>918 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR12</lparam></gate>
<gate>
<ID>764</ID>
<type>DE_TO</type>
<position>137.5,53</position>
<input>
<ID>IN_0</ID>1091 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_LD</lparam></gate>
<gate>
<ID>765</ID>
<type>DE_TO</type>
<position>137.5,47</position>
<input>
<ID>IN_0</ID>1094 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID TR_bus</lparam></gate>
<gate>
<ID>790</ID>
<type>DA_FROM</type>
<position>-118,107.5</position>
<input>
<ID>IN_0</ID>919 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR8</lparam></gate>
<gate>
<ID>275</ID>
<type>DA_FROM</type>
<position>-73,88.5</position>
<input>
<ID>IN_0</ID>324 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR6</lparam></gate>
<gate>
<ID>769</ID>
<type>DE_TO</type>
<position>37,44</position>
<input>
<ID>IN_0</ID>939 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Mem_R</lparam></gate>
<gate>
<ID>781</ID>
<type>DE_TO</type>
<position>-10.5,56.5</position>
<input>
<ID>IN_0</ID>914 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D7</lparam></gate>
<gate>
<ID>785</ID>
<type>DA_FROM</type>
<position>18,48</position>
<input>
<ID>IN_0</ID>922 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D7</lparam></gate>
<gate>
<ID>792</ID>
<type>AA_AND3</type>
<position>24,50</position>
<input>
<ID>IN_0</ID>925 </input>
<input>
<ID>IN_1</ID>923 </input>
<input>
<ID>IN_2</ID>922 </input>
<output>
<ID>OUT</ID>942 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>794</ID>
<type>DA_FROM</type>
<position>18,52</position>
<input>
<ID>IN_0</ID>925 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>800</ID>
<type>AA_AND2</type>
<position>128.5,128</position>
<input>
<ID>IN_0</ID>931 </input>
<input>
<ID>IN_1</ID>992 </input>
<output>
<ID>OUT</ID>930 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>802</ID>
<type>DA_FROM</type>
<position>122,129</position>
<input>
<ID>IN_0</ID>931 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>649</ID>
<type>AA_AND2</type>
<position>24,87.5</position>
<input>
<ID>IN_0</ID>890 </input>
<input>
<ID>IN_1</ID>891 </input>
<output>
<ID>OUT</ID>885 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>806</ID>
<type>DA_FROM</type>
<position>114.5,125.5</position>
<input>
<ID>IN_0</ID>994 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>808</ID>
<type>DA_FROM</type>
<position>114.5,123.5</position>
<input>
<ID>IN_0</ID>993 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>809</ID>
<type>AA_AND2</type>
<position>24,38.5</position>
<input>
<ID>IN_0</ID>935 </input>
<input>
<ID>IN_1</ID>1095 </input>
<output>
<ID>OUT</ID>941 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>810</ID>
<type>DA_FROM</type>
<position>17.5,39.5</position>
<input>
<ID>IN_0</ID>935 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>812</ID>
<type>DA_FROM</type>
<position>10,36.5</position>
<input>
<ID>IN_0</ID>1096 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>813</ID>
<type>DA_FROM</type>
<position>10,34.5</position>
<input>
<ID>IN_0</ID>1097 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>817</ID>
<type>DE_TO</type>
<position>94.5,5</position>
<input>
<ID>IN_0</ID>947 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID SCclr</lparam></gate>
<gate>
<ID>820</ID>
<type>DA_FROM</type>
<position>74,18</position>
<input>
<ID>IN_0</ID>1179 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>821</ID>
<type>DA_FROM</type>
<position>61,23</position>
<input>
<ID>IN_0</ID>1002 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>822</ID>
<type>DA_FROM</type>
<position>61,21</position>
<input>
<ID>IN_0</ID>1001 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1029</ID>
<type>AA_AND2</type>
<position>-83,28.5</position>
<input>
<ID>IN_0</ID>1196 </input>
<input>
<ID>IN_1</ID>1202 </input>
<output>
<ID>OUT</ID>1194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>824</ID>
<type>DE_OR8</type>
<position>87.5,5</position>
<input>
<ID>IN_0</ID>948 </input>
<input>
<ID>IN_1</ID>1178 </input>
<input>
<ID>IN_2</ID>1183 </input>
<input>
<ID>IN_3</ID>1188 </input>
<input>
<ID>IN_4</ID>1062 </input>
<input>
<ID>IN_5</ID>1063 </input>
<input>
<ID>IN_6</ID>1192 </input>
<input>
<ID>IN_7</ID>1191 </input>
<output>
<ID>OUT</ID>947 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>829</ID>
<type>DA_FROM</type>
<position>61,19</position>
<input>
<ID>IN_0</ID>1000 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>836</ID>
<type>AA_AND2</type>
<position>-67,117</position>
<input>
<ID>IN_0</ID>960 </input>
<input>
<ID>IN_1</ID>961 </input>
<output>
<ID>OUT</ID>959 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>838</ID>
<type>DA_FROM</type>
<position>-73,118</position>
<input>
<ID>IN_0</ID>960 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>840</ID>
<type>DA_FROM</type>
<position>-73,116</position>
<input>
<ID>IN_0</ID>961 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>842</ID>
<type>DA_FROM</type>
<position>-73,112.5</position>
<input>
<ID>IN_0</ID>962 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>843</ID>
<type>DA_FROM</type>
<position>-73,110.5</position>
<input>
<ID>IN_0</ID>963 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1024</ID>
<type>AA_AND2</type>
<position>-83,38.5</position>
<input>
<ID>IN_0</ID>1175 </input>
<input>
<ID>IN_1</ID>1176 </input>
<output>
<ID>OUT</ID>1174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>845</ID>
<type>DA_FROM</type>
<position>-129.5,16</position>
<input>
<ID>IN_0</ID>943 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>847</ID>
<type>GA_LED</type>
<position>-59,62</position>
<input>
<ID>N_in2</ID>886 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>868</ID>
<type>AE_OR4</type>
<position>120.5,122.5</position>
<input>
<ID>IN_0</ID>994 </input>
<input>
<ID>IN_1</ID>993 </input>
<input>
<ID>IN_2</ID>995 </input>
<input>
<ID>IN_3</ID>996 </input>
<output>
<ID>OUT</ID>992 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>869</ID>
<type>DA_FROM</type>
<position>114.5,121.5</position>
<input>
<ID>IN_0</ID>995 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>870</ID>
<type>DA_FROM</type>
<position>114.5,119.5</position>
<input>
<ID>IN_0</ID>996 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>871</ID>
<type>AA_AND2</type>
<position>-67,106</position>
<input>
<ID>IN_0</ID>997 </input>
<input>
<ID>IN_1</ID>998 </input>
<output>
<ID>OUT</ID>999 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>873</ID>
<type>DA_FROM</type>
<position>-73,105</position>
<input>
<ID>IN_0</ID>998 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>875</ID>
<type>AE_OR4</type>
<position>67,20</position>
<input>
<ID>IN_0</ID>1002 </input>
<input>
<ID>IN_1</ID>1001 </input>
<input>
<ID>IN_2</ID>1000 </input>
<input>
<ID>IN_3</ID>1004 </input>
<output>
<ID>OUT</ID>1180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>876</ID>
<type>DA_FROM</type>
<position>61,17</position>
<input>
<ID>IN_0</ID>1004 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>48</ID>
<type>DE_TO</type>
<position>22,10</position>
<input>
<ID>IN_0</ID>13 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>926</ID>
<type>DA_FROM</type>
<position>10,32.5</position>
<input>
<ID>IN_0</ID>1098 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>51</ID>
<type>AA_AND3</type>
<position>16,10</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>16 </input>
<input>
<ID>IN_2</ID>15 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>59</ID>
<type>DA_FROM</type>
<position>10,8</position>
<input>
<ID>IN_0</ID>15 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>934</ID>
<type>AA_AND2</type>
<position>65,52.5</position>
<input>
<ID>IN_0</ID>1056 </input>
<input>
<ID>IN_1</ID>1055 </input>
<output>
<ID>OUT</ID>1051 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>10,4</position>
<input>
<ID>IN_0</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D7</lparam></gate>
<gate>
<ID>922</ID>
<type>DA_FROM</type>
<position>72.5,59.5</position>
<input>
<ID>IN_0</ID>1045 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>881</ID>
<type>DA_FROM</type>
<position>-22,92</position>
<input>
<ID>IN_0</ID>1080 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>64</ID>
<type>DE_TO</type>
<position>22,2</position>
<input>
<ID>IN_0</ID>17 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_AND3</type>
<position>16,2</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>20 </input>
<input>
<ID>IN_2</ID>19 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>912</ID>
<type>DA_FROM</type>
<position>72.5,87.5</position>
<input>
<ID>IN_0</ID>1034 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>66</ID>
<type>DA_FROM</type>
<position>10,0</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>885</ID>
<type>AA_AND2</type>
<position>-23,82</position>
<input>
<ID>IN_0</ID>1083 </input>
<input>
<ID>IN_1</ID>1082 </input>
<output>
<ID>OUT</ID>1084 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>DE_TO</type>
<position>-56,55.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /I</lparam></gate>
<gate>
<ID>250</ID>
<type>DE_TO</type>
<position>-61,100.5</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CMA</lparam></gate>
<gate>
<ID>799</ID>
<type>DA_FROM</type>
<position>-126,100.5</position>
<input>
<ID>IN_0</ID>928 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR15</lparam></gate>
<gate>
<ID>972</ID>
<type>AA_AND2</type>
<position>-131,55</position>
<input>
<ID>IN_0</ID>1123 </input>
<input>
<ID>IN_1</ID>1124 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>253</ID>
<type>DA_FROM</type>
<position>-73,101.5</position>
<input>
<ID>IN_0</ID>25 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_AND2</type>
<position>-67,100.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_AND2</type>
<position>-67,95</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>321 </input>
<output>
<ID>OUT</ID>322 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>967</ID>
<type>DA_FROM</type>
<position>-129.5,41.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>265</ID>
<type>DA_FROM</type>
<position>-73,94</position>
<input>
<ID>IN_0</ID>321 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR7</lparam></gate>
<gate>
<ID>269</ID>
<type>DE_TO</type>
<position>-61,89.5</position>
<input>
<ID>IN_0</ID>326 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID CIL</lparam></gate>
<gate>
<ID>271</ID>
<type>DA_FROM</type>
<position>-73,90.5</position>
<input>
<ID>IN_0</ID>323 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>746</ID>
<type>AA_AND2</type>
<position>71.5,128.5</position>
<input>
<ID>IN_0</ID>894 </input>
<input>
<ID>IN_1</ID>895 </input>
<output>
<ID>OUT</ID>893 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>975</ID>
<type>AA_AND2</type>
<position>-123.5,61</position>
<input>
<ID>IN_0</ID>1125 </input>
<input>
<ID>IN_1</ID>1126 </input>
<output>
<ID>OUT</ID>1127 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>273</ID>
<type>AA_AND2</type>
<position>-67,89.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>324 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>DE_TO</type>
<position>-61,84</position>
<input>
<ID>IN_0</ID>350 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID INP</lparam></gate>
<gate>
<ID>963</ID>
<type>DA_FROM</type>
<position>66,112</position>
<input>
<ID>IN_0</ID>957 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND2</type>
<position>-67,84</position>
<input>
<ID>IN_0</ID>337 </input>
<input>
<ID>IN_1</ID>349 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>983</ID>
<type>DA_FROM</type>
<position>132.5,34</position>
<input>
<ID>IN_0</ID>1058 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>991</ID>
<type>AE_SMALL_INVERTER</type>
<position>-89,-0.5</position>
<input>
<ID>IN_0</ID>1162 </input>
<output>
<ID>OUT_0</ID>1172 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>289</ID>
<type>BE_JKFF_LOW</type>
<position>-116.5,1.5</position>
<input>
<ID>J</ID>1140 </input>
<input>
<ID>K</ID>83 </input>
<output>
<ID>Q</ID>417 </output>
<input>
<ID>clock</ID>352 </input>
<output>
<ID>nQ</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>291</ID>
<type>DE_TO</type>
<position>-109.5,3.5</position>
<input>
<ID>IN_0</ID>417 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>293</ID>
<type>GA_LED</type>
<position>-112.5,6</position>
<input>
<ID>N_in2</ID>417 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>979</ID>
<type>DA_FROM</type>
<position>132.5,90.5</position>
<input>
<ID>IN_0</ID>1057 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>295</ID>
<type>DE_TO</type>
<position>-51,24</position>
<input>
<ID>IN_0</ID>418 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /E</lparam></gate>
<gate>
<ID>999</ID>
<type>DE_TO</type>
<position>-9.5,11</position>
<input>
<ID>IN_0</ID>1138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /T1</lparam></gate>
<gate>
<ID>297</ID>
<type>BE_JKFF_LOW</type>
<position>-58,26</position>
<input>
<ID>J</ID>1153 </input>
<input>
<ID>K</ID>1060 </input>
<output>
<ID>Q</ID>444 </output>
<input>
<ID>clock</ID>443 </input>
<output>
<ID>nQ</ID>418 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>992</ID>
<type>DA_FROM</type>
<position>-94,-0.5</position>
<input>
<ID>IN_0</ID>1162 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>145</ID>
<type>AE_OR2</type>
<position>131,99</position>
<input>
<ID>IN_0</ID>884 </input>
<input>
<ID>IN_1</ID>786 </input>
<output>
<ID>OUT</ID>1009 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>298</ID>
<type>DE_TO</type>
<position>-51,28</position>
<input>
<ID>IN_0</ID>444 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>299</ID>
<type>GA_LED</type>
<position>-54,30.5</position>
<input>
<ID>N_in2</ID>444 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>301</ID>
<type>DA_FROM</type>
<position>-122.5,57.5</position>
<input>
<ID>IN_0</ID>470 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>987</ID>
<type>DA_FROM</type>
<position>-22,86</position>
<input>
<ID>IN_0</ID>1129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>1007</ID>
<type>DA_FROM</type>
<position>-135.5,4.5</position>
<input>
<ID>IN_0</ID>1144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /T2</lparam></gate>
<gate>
<ID>512</ID>
<type>DA_FROM</type>
<position>125.5,70</position>
<input>
<ID>IN_0</ID>1014 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>305</ID>
<type>DA_FROM</type>
<position>-122.5,31.5</position>
<input>
<ID>IN_0</ID>713 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>307</ID>
<type>DA_FROM</type>
<position>-122.5,44</position>
<input>
<ID>IN_0</ID>688 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>995</ID>
<type>AE_SMALL_INVERTER</type>
<position>-13,13</position>
<input>
<ID>IN_0</ID>411 </input>
<output>
<ID>OUT_0</ID>1137 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>309</ID>
<type>DE_TO</type>
<position>-109.5,55.5</position>
<input>
<ID>IN_0</ID>469 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /IEN</lparam></gate>
<gate>
<ID>311</ID>
<type>BE_JKFF_LOW</type>
<position>-116.5,44</position>
<input>
<ID>J</ID>1116 </input>
<input>
<ID>K</ID>1118 </input>
<output>
<ID>Q</ID>707 </output>
<input>
<ID>clock</ID>688 </input>
<output>
<ID>nQ</ID>687 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>1015</ID>
<type>AE_OR2</type>
<position>-143.5,4.5</position>
<input>
<ID>IN_0</ID>1151 </input>
<input>
<ID>IN_1</ID>1150 </input>
<output>
<ID>OUT</ID>1149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>313</ID>
<type>DE_TO</type>
<position>-109.5,46</position>
<input>
<ID>IN_0</ID>707 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>1008</ID>
<type>DA_FROM</type>
<position>-135.5,2.5</position>
<input>
<ID>IN_0</ID>1145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /T1</lparam></gate>
<gate>
<ID>314</ID>
<type>GA_LED</type>
<position>-112.5,48.5</position>
<input>
<ID>N_in2</ID>707 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>315</ID>
<type>DE_TO</type>
<position>-109.5,29.5</position>
<input>
<ID>IN_0</ID>709 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /FGO</lparam></gate>
<gate>
<ID>319</ID>
<type>BE_JKFF_LOW</type>
<position>-116.5,31.5</position>
<input>
<ID>J</ID>1115 </input>
<input>
<ID>K</ID>1117 </input>
<output>
<ID>Q</ID>714 </output>
<input>
<ID>clock</ID>713 </input>
<output>
<ID>nQ</ID>709 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>322</ID>
<type>DE_TO</type>
<position>-109.5,33.5</position>
<input>
<ID>IN_0</ID>714 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>349</ID>
<type>GA_LED</type>
<position>-112.5,36</position>
<input>
<ID>N_in2</ID>714 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>403</ID>
<type>AE_OR2</type>
<position>16.5,128.5</position>
<input>
<ID>IN_0</ID>759 </input>
<input>
<ID>IN_1</ID>760 </input>
<output>
<ID>OUT</ID>734 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>430</ID>
<type>AE_OR2</type>
<position>31,124</position>
<input>
<ID>IN_0</ID>739 </input>
<input>
<ID>IN_1</ID>761 </input>
<output>
<ID>OUT</ID>735 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>457</ID>
<type>DA_FROM</type>
<position>18,125</position>
<input>
<ID>IN_0</ID>740 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>814</ID>
<type>AE_OR3</type>
<position>-29,122.5</position>
<input>
<ID>IN_0</ID>1076 </input>
<input>
<ID>IN_1</ID>1077 </input>
<input>
<ID>IN_2</ID>1075 </input>
<output>
<ID>OUT</ID>1074 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>484</ID>
<type>DA_FROM</type>
<position>10.5,129.5</position>
<input>
<ID>IN_0</ID>759 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>511</ID>
<type>DA_FROM</type>
<position>10.5,127.5</position>
<input>
<ID>IN_0</ID>760 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>513</ID>
<type>AA_AND3</type>
<position>24,120</position>
<input>
<ID>IN_0</ID>765 </input>
<input>
<ID>IN_1</ID>766 </input>
<input>
<ID>IN_2</ID>785 </input>
<output>
<ID>OUT</ID>761 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>519</ID>
<type>DA_FROM</type>
<position>18,122</position>
<input>
<ID>IN_0</ID>765 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /D7</lparam></gate>
<gate>
<ID>521</ID>
<type>DA_FROM</type>
<position>18,120</position>
<input>
<ID>IN_0</ID>766 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID I</lparam></gate>
<gate>
<ID>525</ID>
<type>DA_FROM</type>
<position>18,118</position>
<input>
<ID>IN_0</ID>785 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T3</lparam></gate>
<gate>
<ID>548</ID>
<type>AA_AND2</type>
<position>24,106</position>
<input>
<ID>IN_0</ID>787 </input>
<input>
<ID>IN_1</ID>791 </input>
<output>
<ID>OUT</ID>955 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>899</ID>
<type>AA_AND3</type>
<position>78.5,85.5</position>
<input>
<ID>IN_0</ID>1034 </input>
<input>
<ID>IN_1</ID>1036 </input>
<input>
<ID>IN_2</ID>1048 </input>
<output>
<ID>OUT</ID>1023 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>552</ID>
<type>DA_FROM</type>
<position>18,107</position>
<input>
<ID>IN_0</ID>787 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>919</ID>
<type>DA_FROM</type>
<position>72.5,76.5</position>
<input>
<ID>IN_0</ID>1042 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>1069</ID>
<type>DA_FROM</type>
<position>74,1.5</position>
<input>
<ID>IN_0</ID>1191 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>591</ID>
<type>DA_FROM</type>
<position>25,99</position>
<input>
<ID>IN_0</ID>881 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>595</ID>
<type>AA_AND2</type>
<position>31,100</position>
<input>
<ID>IN_0</ID>880 </input>
<input>
<ID>IN_1</ID>881 </input>
<output>
<ID>OUT</ID>882 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>617</ID>
<type>DA_FROM</type>
<position>25,101</position>
<input>
<ID>IN_0</ID>880 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>619</ID>
<type>AE_OR2</type>
<position>31,89.5</position>
<input>
<ID>IN_0</ID>887 </input>
<input>
<ID>IN_1</ID>885 </input>
<output>
<ID>OUT</ID>883 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>645</ID>
<type>AA_AND2</type>
<position>24,91.5</position>
<input>
<ID>IN_0</ID>888 </input>
<input>
<ID>IN_1</ID>889 </input>
<output>
<ID>OUT</ID>887 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>798</ID>
<type>DA_FROM</type>
<position>-118,101.5</position>
<input>
<ID>IN_0</ID>920 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR14</lparam></gate>
<gate>
<ID>1030</ID>
<type>DA_FROM</type>
<position>-89,34.5</position>
<input>
<ID>IN_0</ID>1195 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR7</lparam></gate>
<gate>
<ID>672</ID>
<type>DA_FROM</type>
<position>18,92.5</position>
<input>
<ID>IN_0</ID>888 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>676</ID>
<type>DA_FROM</type>
<position>18,90.5</position>
<input>
<ID>IN_0</ID>889 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>884</ID>
<type>DA_FROM</type>
<position>-29,83</position>
<input>
<ID>IN_0</ID>1083 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>723</ID>
<type>DA_FROM</type>
<position>18,88.5</position>
<input>
<ID>IN_0</ID>890 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>772</ID>
<type>DA_FROM</type>
<position>-28,101.5</position>
<input>
<ID>IN_0</ID>1072 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>739</ID>
<type>DA_FROM</type>
<position>18,86.5</position>
<input>
<ID>IN_0</ID>891 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>741</ID>
<type>AA_AND2</type>
<position>71.5,124.5</position>
<input>
<ID>IN_0</ID>896 </input>
<input>
<ID>IN_1</ID>897 </input>
<output>
<ID>OUT</ID>892 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>894</ID>
<type>AA_AND2</type>
<position>78.5,103.5</position>
<input>
<ID>IN_0</ID>1027 </input>
<input>
<ID>IN_1</ID>1028 </input>
<output>
<ID>OUT</ID>1026 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>888</ID>
<type>AA_AND2</type>
<position>-16,77</position>
<input>
<ID>IN_0</ID>1086 </input>
<input>
<ID>IN_1</ID>1085 </input>
<output>
<ID>OUT</ID>1087 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>743</ID>
<type>AE_OR2</type>
<position>78.5,126.5</position>
<input>
<ID>IN_0</ID>893 </input>
<input>
<ID>IN_1</ID>892 </input>
<output>
<ID>OUT</ID>900 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>DA_FROM</type>
<position>118,98</position>
<input>
<ID>IN_0</ID>901 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>747</ID>
<type>DA_FROM</type>
<position>65.5,129.5</position>
<input>
<ID>IN_0</ID>894 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D4</lparam></gate>
<gate>
<ID>780</ID>
<type>DA_FROM</type>
<position>-126,114.5</position>
<input>
<ID>IN_0</ID>924 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR1</lparam></gate>
<gate>
<ID>749</ID>
<type>DA_FROM</type>
<position>65.5,127.5</position>
<input>
<ID>IN_0</ID>895 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>774</ID>
<type>DE_OR8</type>
<position>-112,104</position>
<input>
<ID>IN_0</ID>919 </input>
<input>
<ID>IN_1</ID>929 </input>
<input>
<ID>IN_2</ID>917 </input>
<input>
<ID>IN_3</ID>933 </input>
<input>
<ID>IN_4</ID>928 </input>
<input>
<ID>IN_5</ID>920 </input>
<input>
<ID>IN_6</ID>932 </input>
<input>
<ID>IN_7</ID>918 </input>
<output>
<ID>OUT</ID>911 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>753</ID>
<type>DA_FROM</type>
<position>65.5,123.5</position>
<input>
<ID>IN_0</ID>897 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>778</ID>
<type>DA_FROM</type>
<position>-118,115.5</position>
<input>
<ID>IN_0</ID>912 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR0</lparam></gate>
<gate>
<ID>755</ID>
<type>AE_OR3</type>
<position>-65,21.5</position>
<input>
<ID>IN_0</ID>1061 </input>
<input>
<ID>IN_1</ID>1142 </input>
<input>
<ID>IN_2</ID>1148 </input>
<output>
<ID>OUT</ID>1060 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>788</ID>
<type>DA_FROM</type>
<position>-118,109.5</position>
<input>
<ID>IN_0</ID>915 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR6</lparam></gate>
<gate>
<ID>757</ID>
<type>AA_AND2</type>
<position>-72.5,16.5</position>
<input>
<ID>IN_0</ID>1143 </input>
<input>
<ID>IN_1</ID>1147 </input>
<output>
<ID>OUT</ID>1142 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>782</ID>
<type>DA_FROM</type>
<position>-118,113.5</position>
<input>
<ID>IN_0</ID>916 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR2</lparam></gate>
<gate>
<ID>767</ID>
<type>DA_FROM</type>
<position>-28,99.5</position>
<input>
<ID>IN_0</ID>1071 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR11</lparam></gate>
<gate>
<ID>784</ID>
<type>DA_FROM</type>
<position>-126,112.5</position>
<input>
<ID>IN_0</ID>926 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR3</lparam></gate>
<gate>
<ID>787</ID>
<type>DA_FROM</type>
<position>-126,110.5</position>
<input>
<ID>IN_0</ID>927 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR5</lparam></gate>
<gate>
<ID>789</ID>
<type>DA_FROM</type>
<position>-126,108.5</position>
<input>
<ID>IN_0</ID>921 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR7</lparam></gate>
<gate>
<ID>793</ID>
<type>DA_FROM</type>
<position>-118,105.5</position>
<input>
<ID>IN_0</ID>917 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR10</lparam></gate>
<gate>
<ID>795</ID>
<type>DA_FROM</type>
<position>-126,104.5</position>
<input>
<ID>IN_0</ID>933 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR11</lparam></gate>
<gate>
<ID>797</ID>
<type>DA_FROM</type>
<position>-126,102.5</position>
<input>
<ID>IN_0</ID>932 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR13</lparam></gate>
<gate>
<ID>804</ID>
<type>BE_NOR2</type>
<position>-104,89</position>
<input>
<ID>IN_0</ID>944 </input>
<input>
<ID>IN_1</ID>945 </input>
<output>
<ID>OUT</ID>1007 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>805</ID>
<type>DE_OR8</type>
<position>-112,93</position>
<input>
<ID>IN_0</ID>965 </input>
<input>
<ID>IN_1</ID>983 </input>
<input>
<ID>IN_2</ID>967 </input>
<input>
<ID>IN_3</ID>982 </input>
<input>
<ID>IN_4</ID>1006 </input>
<input>
<ID>IN_5</ID>977 </input>
<input>
<ID>IN_6</ID>1005 </input>
<input>
<ID>IN_7</ID>976 </input>
<output>
<ID>OUT</ID>944 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>807</ID>
<type>DE_OR8</type>
<position>-112,85</position>
<input>
<ID>IN_0</ID>951 </input>
<input>
<ID>IN_1</ID>981 </input>
<input>
<ID>IN_2</ID>952 </input>
<input>
<ID>IN_3</ID>980 </input>
<input>
<ID>IN_4</ID>979 </input>
<input>
<ID>IN_5</ID>953 </input>
<input>
<ID>IN_6</ID>978 </input>
<input>
<ID>IN_7</ID>950 </input>
<output>
<ID>OUT</ID>945 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>671</ID>
<type>AA_AND2</type>
<position>-83,10.5</position>
<input>
<ID>IN_0</ID>938 </input>
<input>
<ID>IN_1</ID>1010 </input>
<output>
<ID>OUT</ID>908 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>816</ID>
<type>DA_FROM</type>
<position>-118,96.5</position>
<input>
<ID>IN_0</ID>965 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>818</ID>
<type>DA_FROM</type>
<position>-127.5,95.5</position>
<input>
<ID>IN_0</ID>983 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo1</lparam></gate>
<gate>
<ID>825</ID>
<type>DA_FROM</type>
<position>-127.5,93.5</position>
<input>
<ID>IN_0</ID>982 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo3</lparam></gate>
<gate>
<ID>1034</ID>
<type>DA_FROM</type>
<position>-89,32.5</position>
<input>
<ID>IN_0</ID>1203 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>827</ID>
<type>DA_FROM</type>
<position>-118,92.5</position>
<input>
<ID>IN_0</ID>976 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo4</lparam></gate>
<gate>
<ID>828</ID>
<type>DA_FROM</type>
<position>-127.5,91.5</position>
<input>
<ID>IN_0</ID>1005 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo5</lparam></gate>
<gate>
<ID>835</ID>
<type>DA_FROM</type>
<position>-118,90.5</position>
<input>
<ID>IN_0</ID>977 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo6</lparam></gate>
<gate>
<ID>839</ID>
<type>DA_FROM</type>
<position>-118,88.5</position>
<input>
<ID>IN_0</ID>951 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo8</lparam></gate>
<gate>
<ID>844</ID>
<type>DA_FROM</type>
<position>-127.5,87.5</position>
<input>
<ID>IN_0</ID>981 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo9</lparam></gate>
<gate>
<ID>846</ID>
<type>DA_FROM</type>
<position>-118,86.5</position>
<input>
<ID>IN_0</ID>952 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo10</lparam></gate>
<gate>
<ID>848</ID>
<type>DA_FROM</type>
<position>-127.5,85.5</position>
<input>
<ID>IN_0</ID>980 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo11</lparam></gate>
<gate>
<ID>1</ID>
<type>AA_AND2</type>
<position>-123.5,-3</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>850</ID>
<type>DA_FROM</type>
<position>-127.5,83.5</position>
<input>
<ID>IN_0</ID>978 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo13</lparam></gate>
<gate>
<ID>1027</ID>
<type>AA_LABEL</type>
<position>26.5,133.5</position>
<gparam>LABEL_TEXT AR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>867</ID>
<type>DA_FROM</type>
<position>-118,82.5</position>
<input>
<ID>IN_0</ID>953 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo14</lparam></gate>
<gate>
<ID>874</ID>
<type>DA_FROM</type>
<position>-127.5,81.5</position>
<input>
<ID>IN_0</ID>979 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>878</ID>
<type>DE_TO</type>
<position>-98,89</position>
<input>
<ID>IN_0</ID>1007 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID AC=0</lparam></gate>
<gate>
<ID>896</ID>
<type>AA_AND2</type>
<position>78.5,98.5</position>
<input>
<ID>IN_0</ID>1030 </input>
<input>
<ID>IN_1</ID>1029 </input>
<output>
<ID>OUT</ID>1025 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>898</ID>
<type>AA_AND3</type>
<position>78.5,92.5</position>
<input>
<ID>IN_0</ID>1031 </input>
<input>
<ID>IN_1</ID>1033 </input>
<input>
<ID>IN_2</ID>1032 </input>
<output>
<ID>OUT</ID>1024 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>900</ID>
<type>AA_AND3</type>
<position>78.5,78.5</position>
<input>
<ID>IN_0</ID>1041 </input>
<input>
<ID>IN_1</ID>1043 </input>
<input>
<ID>IN_2</ID>1042 </input>
<output>
<ID>OUT</ID>1022 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1049</ID>
<type>AA_LABEL</type>
<position>77,27.5</position>
<gparam>LABEL_TEXT Sequence Counter Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>901</ID>
<type>AA_AND3</type>
<position>78.5,71.5</position>
<input>
<ID>IN_0</ID>1038 </input>
<input>
<ID>IN_1</ID>1037 </input>
<input>
<ID>IN_2</ID>1039 </input>
<output>
<ID>OUT</ID>1021 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>902</ID>
<type>AA_AND3</type>
<position>78.5,64.5</position>
<input>
<ID>IN_0</ID>1040 </input>
<input>
<ID>IN_1</ID>1047 </input>
<input>
<ID>IN_2</ID>1046 </input>
<output>
<ID>OUT</ID>1020 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>904</ID>
<type>AA_AND2</type>
<position>78.5,58.5</position>
<input>
<ID>IN_0</ID>1045 </input>
<input>
<ID>IN_1</ID>1050 </input>
<output>
<ID>OUT</ID>1019 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>905</ID>
<type>DA_FROM</type>
<position>72.5,102.5</position>
<input>
<ID>IN_0</ID>1028 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>906</ID>
<type>DA_FROM</type>
<position>72.5,104.5</position>
<input>
<ID>IN_0</ID>1027 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>907</ID>
<type>DA_FROM</type>
<position>72.5,97.5</position>
<input>
<ID>IN_0</ID>1029 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>908</ID>
<type>DA_FROM</type>
<position>72.5,99.5</position>
<input>
<ID>IN_0</ID>1030 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1057</ID>
<type>AA_LABEL</type>
<position>131,133.5</position>
<gparam>LABEL_TEXT DR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>909</ID>
<type>DA_FROM</type>
<position>72.5,94.5</position>
<input>
<ID>IN_0</ID>1031 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>910</ID>
<type>DA_FROM</type>
<position>72.5,90.5</position>
<input>
<ID>IN_0</ID>1032 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR=0</lparam></gate>
<gate>
<ID>911</ID>
<type>DA_FROM</type>
<position>72.5,92.5</position>
<input>
<ID>IN_0</ID>1033 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>914</ID>
<type>DA_FROM</type>
<position>72.5,85.5</position>
<input>
<ID>IN_0</ID>1036 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR4</lparam></gate>
<gate>
<ID>915</ID>
<type>DA_FROM</type>
<position>72.5,71.5</position>
<input>
<ID>IN_0</ID>1037 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR2</lparam></gate>
<gate>
<ID>1065</ID>
<type>AA_AND2</type>
<position>80,5.5</position>
<input>
<ID>IN_0</ID>1190 </input>
<input>
<ID>IN_1</ID>1189 </input>
<output>
<ID>OUT</ID>1188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_AND2</type>
<position>124,97</position>
<input>
<ID>IN_0</ID>901 </input>
<input>
<ID>IN_1</ID>946 </input>
<output>
<ID>OUT</ID>786 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>916</ID>
<type>DA_FROM</type>
<position>72.5,80.5</position>
<input>
<ID>IN_0</ID>1041 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>918</ID>
<type>DA_FROM</type>
<position>72.5,73.5</position>
<input>
<ID>IN_0</ID>1038 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>920</ID>
<type>DA_FROM</type>
<position>72.5,66.5</position>
<input>
<ID>IN_0</ID>1040 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>923</ID>
<type>DA_FROM</type>
<position>72.5,62.5</position>
<input>
<ID>IN_0</ID>1046 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /E</lparam></gate>
<gate>
<ID>924</ID>
<type>DA_FROM</type>
<position>72.5,64.5</position>
<input>
<ID>IN_0</ID>1047 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR1</lparam></gate>
<gate>
<ID>1073</ID>
<type>DA_FROM</type>
<position>74,-4.5</position>
<input>
<ID>IN_0</ID>1063 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>927</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,83.5</position>
<input>
<ID>IN_0</ID>1049 </input>
<output>
<ID>OUT_0</ID>1048 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>929</ID>
<type>DA_FROM</type>
<position>67.5,83.5</position>
<input>
<ID>IN_0</ID>1049 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>931</ID>
<type>AE_OR2</type>
<position>71.5,55</position>
<input>
<ID>IN_0</ID>1052 </input>
<input>
<ID>IN_1</ID>1051 </input>
<output>
<ID>OUT</ID>1050 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>935</ID>
<type>DA_FROM</type>
<position>59,58.5</position>
<input>
<ID>IN_0</ID>1054 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR8</lparam></gate>
<gate>
<ID>936</ID>
<type>DA_FROM</type>
<position>59,56.5</position>
<input>
<ID>IN_0</ID>1053 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>937</ID>
<type>DA_FROM</type>
<position>59,53.5</position>
<input>
<ID>IN_0</ID>1056 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR9</lparam></gate>
<gate>
<ID>938</ID>
<type>DA_FROM</type>
<position>59,51.5</position>
<input>
<ID>IN_0</ID>1055 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>944</ID>
<type>AA_AND2</type>
<position>72,42.5</position>
<input>
<ID>IN_0</ID>1066 </input>
<input>
<ID>IN_1</ID>1065 </input>
<output>
<ID>OUT</ID>1069 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>948</ID>
<type>DA_FROM</type>
<position>72,46.5</position>
<input>
<ID>IN_0</ID>1068 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>949</ID>
<type>DA_FROM</type>
<position>66,43.5</position>
<input>
<ID>IN_0</ID>1066 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>950</ID>
<type>DA_FROM</type>
<position>66,41.5</position>
<input>
<ID>IN_0</ID>1065 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>952</ID>
<type>AE_OR2</type>
<position>78.5,44.5</position>
<input>
<ID>IN_0</ID>1068 </input>
<input>
<ID>IN_1</ID>1069 </input>
<output>
<ID>OUT</ID>1067 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_AND2</type>
<position>131.5,110.5</position>
<input>
<ID>IN_0</ID>413 </input>
<input>
<ID>IN_1</ID>681 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>DA_FROM</type>
<position>125.5,111.5</position>
<input>
<ID>IN_0</ID>413 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>60</ID>
<type>DA_FROM</type>
<position>125.5,109.5</position>
<input>
<ID>IN_0</ID>681 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_AND2</type>
<position>124,101</position>
<input>
<ID>IN_0</ID>898 </input>
<input>
<ID>IN_1</ID>899 </input>
<output>
<ID>OUT</ID>884 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>971</ID>
<type>DA_FROM</type>
<position>-137,56</position>
<input>
<ID>IN_0</ID>1123 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>285</ID>
<type>DA_FROM</type>
<position>118,100</position>
<input>
<ID>IN_0</ID>899 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>300</ID>
<type>DA_FROM</type>
<position>118,96</position>
<input>
<ID>IN_0</ID>946 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>377</ID>
<type>AA_AND4</type>
<position>-72.5,9.5</position>
<input>
<ID>IN_0</ID>904 </input>
<input>
<ID>IN_1</ID>908 </input>
<input>
<ID>IN_2</ID>1154 </input>
<input>
<ID>IN_3</ID>1157 </input>
<output>
<ID>OUT</ID>1148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1070</ID>
<type>DA_FROM</type>
<position>74,-1.5</position>
<input>
<ID>IN_0</ID>1192 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>697</ID>
<type>DE_TO</type>
<position>137.5,90.5</position>
<input>
<ID>IN_0</ID>1057 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID DR_CLR</lparam></gate>
<gate>
<ID>404</ID>
<type>AA_AND2</type>
<position>131.5,74.5</position>
<input>
<ID>IN_0</ID>1011 </input>
<input>
<ID>IN_1</ID>1012 </input>
<output>
<ID>OUT</ID>1013 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>431</ID>
<type>DA_FROM</type>
<position>125.5,75.5</position>
<input>
<ID>IN_0</ID>1011 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>623</ID>
<type>AA_AND2</type>
<position>-22,113</position>
<input>
<ID>IN_0</ID>1044 </input>
<input>
<ID>IN_1</ID>906 </input>
<output>
<ID>OUT</ID>1018 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>458</ID>
<type>DA_FROM</type>
<position>125.5,73.5</position>
<input>
<ID>IN_0</ID>1012 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>485</ID>
<type>AA_AND2</type>
<position>131.5,69</position>
<input>
<ID>IN_0</ID>1014 </input>
<input>
<ID>IN_1</ID>1015 </input>
<output>
<ID>OUT</ID>1016 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>515</ID>
<type>DA_FROM</type>
<position>125.5,68</position>
<input>
<ID>IN_0</ID>1015 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>549</ID>
<type>AE_OR3</type>
<position>-15,113</position>
<input>
<ID>IN_0</ID>1073 </input>
<input>
<ID>IN_1</ID>1018 </input>
<input>
<ID>IN_2</ID>1070 </input>
<output>
<ID>OUT</ID>1017 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1054</ID>
<type>DA_FROM</type>
<position>74,13.5</position>
<input>
<ID>IN_0</ID>1182 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>696</ID>
<type>DA_FROM</type>
<position>-28,114</position>
<input>
<ID>IN_0</ID>1044 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID r</lparam></gate>
<gate>
<ID>724</ID>
<type>DA_FROM</type>
<position>-35,111.5</position>
<input>
<ID>IN_0</ID>905 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR9</lparam></gate>
<gate>
<ID>886</ID>
<type>DA_FROM</type>
<position>-22,76</position>
<input>
<ID>IN_0</ID>1085 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>733</ID>
<type>DA_FROM</type>
<position>-35,109.5</position>
<input>
<ID>IN_0</ID>902 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR7</lparam></gate>
<gate>
<ID>777</ID>
<type>AA_AND2</type>
<position>-22,119</position>
<input>
<ID>IN_0</ID>1074 </input>
<input>
<ID>IN_1</ID>1078 </input>
<output>
<ID>OUT</ID>1073 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>830</ID>
<type>DA_FROM</type>
<position>-35,120.5</position>
<input>
<ID>IN_0</ID>1075 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>831</ID>
<type>DA_FROM</type>
<position>-35,124.5</position>
<input>
<ID>IN_0</ID>1076 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D0</lparam></gate>
<gate>
<ID>832</ID>
<type>DA_FROM</type>
<position>-35,122.5</position>
<input>
<ID>IN_0</ID>1077 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>879</ID>
<type>AA_AND2</type>
<position>-16,91</position>
<input>
<ID>IN_0</ID>1080 </input>
<input>
<ID>IN_1</ID>1079 </input>
<output>
<ID>OUT</ID>1064 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>883</ID>
<type>DA_FROM</type>
<position>-29,81</position>
<input>
<ID>IN_0</ID>1082 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR11</lparam></gate>
<gate>
<ID>887</ID>
<type>DA_FROM</type>
<position>-22,78</position>
<input>
<ID>IN_0</ID>1086 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>1072</ID>
<type>FF_GND</type>
<position>84,-5.5</position>
<output>
<ID>OUT_0</ID>1062 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>893</ID>
<type>DA_FROM</type>
<position>125.5,52</position>
<input>
<ID>IN_0</ID>1090 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T0</lparam></gate>
<gate>
<ID>895</ID>
<type>DA_FROM</type>
<position>125.5,48</position>
<input>
<ID>IN_0</ID>1092 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>897</ID>
<type>AA_AND2</type>
<position>131.5,47</position>
<input>
<ID>IN_0</ID>1092 </input>
<input>
<ID>IN_1</ID>1093 </input>
<output>
<ID>OUT</ID>1094 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>903</ID>
<type>DA_FROM</type>
<position>125.5,46</position>
<input>
<ID>IN_0</ID>1093 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>928</ID>
<type>DA_FROM</type>
<position>10,30.5</position>
<input>
<ID>IN_0</ID>1099 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>932</ID>
<type>AA_AND2</type>
<position>24,44</position>
<input>
<ID>IN_0</ID>1102 </input>
<input>
<ID>IN_1</ID>1101 </input>
<output>
<ID>OUT</ID>1100 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>939</ID>
<type>DA_FROM</type>
<position>18,45</position>
<input>
<ID>IN_0</ID>1102 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /R</lparam></gate>
<gate>
<ID>941</ID>
<type>AE_OR3</type>
<position>31,66</position>
<input>
<ID>IN_0</ID>1106 </input>
<input>
<ID>IN_1</ID>1104 </input>
<input>
<ID>IN_2</ID>1105 </input>
<output>
<ID>OUT</ID>1103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>943</ID>
<type>AA_AND2</type>
<position>24,66</position>
<input>
<ID>IN_0</ID>1110 </input>
<input>
<ID>IN_1</ID>1107 </input>
<output>
<ID>OUT</ID>1104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>945</ID>
<type>AA_AND2</type>
<position>24,71</position>
<input>
<ID>IN_0</ID>1108 </input>
<input>
<ID>IN_1</ID>1109 </input>
<output>
<ID>OUT</ID>1106 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>946</ID>
<type>AA_AND2</type>
<position>24,57.5</position>
<input>
<ID>IN_0</ID>1113 </input>
<input>
<ID>IN_1</ID>1114 </input>
<output>
<ID>OUT</ID>1105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>951</ID>
<type>AE_OR2</type>
<position>17,62.5</position>
<input>
<ID>IN_0</ID>1111 </input>
<input>
<ID>IN_1</ID>1112 </input>
<output>
<ID>OUT</ID>1107 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>DE_TO</type>
<position>139,18</position>
<input>
<ID>IN_0</ID>85 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID OUTR_LD</lparam></gate>
<gate>
<ID>953</ID>
<type>DA_FROM</type>
<position>18,72</position>
<input>
<ID>IN_0</ID>1108 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>954</ID>
<type>DA_FROM</type>
<position>18,70</position>
<input>
<ID>IN_0</ID>1109 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>955</ID>
<type>DA_FROM</type>
<position>18,67</position>
<input>
<ID>IN_0</ID>1110 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>956</ID>
<type>DA_FROM</type>
<position>11,63.5</position>
<input>
<ID>IN_0</ID>1111 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>957</ID>
<type>DA_FROM</type>
<position>11,61.5</position>
<input>
<ID>IN_0</ID>1112 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D5</lparam></gate>
<gate>
<ID>958</ID>
<type>DA_FROM</type>
<position>18,58.5</position>
<input>
<ID>IN_0</ID>1113 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>959</ID>
<type>DA_FROM</type>
<position>18,56.5</position>
<input>
<ID>IN_0</ID>1114 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D6</lparam></gate>
<gate>
<ID>961</ID>
<type>DA_FROM</type>
<position>-122.5,33.5</position>
<input>
<ID>IN_0</ID>1115 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO_SET</lparam></gate>
<gate>
<ID>962</ID>
<type>DA_FROM</type>
<position>-122.5,46</position>
<input>
<ID>IN_0</ID>1116 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI_SET</lparam></gate>
<gate>
<ID>964</ID>
<type>AA_AND2</type>
<position>-123.5,28</position>
<input>
<ID>IN_0</ID>1121 </input>
<input>
<ID>IN_1</ID>1122 </input>
<output>
<ID>OUT</ID>1117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>965</ID>
<type>AA_AND2</type>
<position>-123.5,40.5</position>
<input>
<ID>IN_0</ID>1119 </input>
<input>
<ID>IN_1</ID>1120 </input>
<output>
<ID>OUT</ID>1118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>968</ID>
<type>DA_FROM</type>
<position>-129.5,39.5</position>
<input>
<ID>IN_0</ID>1120 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR11</lparam></gate>
<gate>
<ID>969</ID>
<type>DA_FROM</type>
<position>-129.5,29</position>
<input>
<ID>IN_0</ID>1121 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>970</ID>
<type>DA_FROM</type>
<position>-129.5,27</position>
<input>
<ID>IN_0</ID>1122 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR10</lparam></gate>
<gate>
<ID>973</ID>
<type>DA_FROM</type>
<position>-137,54</position>
<input>
<ID>IN_0</ID>1124 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR6</lparam></gate>
<gate>
<ID>974</ID>
<type>DA_FROM</type>
<position>-129.5,62</position>
<input>
<ID>IN_0</ID>1125 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>976</ID>
<type>DA_FROM</type>
<position>-129.5,60</position>
<input>
<ID>IN_0</ID>1126 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR7</lparam></gate>
<gate>
<ID>980</ID>
<type>AA_AND2</type>
<position>-80,57.5</position>
<input>
<ID>IN_0</ID>1135 </input>
<input>
<ID>IN_1</ID>1136 </input>
<output>
<ID>OUT</ID>1134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>982</ID>
<type>AA_AND2</type>
<position>-70,61</position>
<input>
<ID>IN_0</ID>1132 </input>
<input>
<ID>IN_1</ID>1134 </input>
<output>
<ID>OUT</ID>1130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>984</ID>
<type>AA_AND2</type>
<position>-70,54</position>
<input>
<ID>IN_0</ID>1133 </input>
<input>
<ID>IN_1</ID>1134 </input>
<output>
<ID>OUT</ID>1131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>986</ID>
<type>AE_SMALL_INVERTER</type>
<position>-75,57.5</position>
<input>
<ID>IN_0</ID>1132 </input>
<output>
<ID>OUT_0</ID>1133 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>989</ID>
<type>DA_FROM</type>
<position>-86,56.5</position>
<input>
<ID>IN_0</ID>1136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>997</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16,9</position>
<input>
<ID>IN_0</ID>406 </input>
<output>
<ID>OUT_0</ID>1139 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>998</ID>
<type>DE_TO</type>
<position>-8,13</position>
<input>
<ID>IN_0</ID>1137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /T0</lparam></gate>
<gate>
<ID>1002</ID>
<type>AA_AND4</type>
<position>-129.5,3.5</position>
<input>
<ID>IN_0</ID>1141 </input>
<input>
<ID>IN_1</ID>1144 </input>
<input>
<ID>IN_2</ID>1145 </input>
<input>
<ID>IN_3</ID>1146 </input>
<output>
<ID>OUT</ID>1140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>1025</ID>
<type>AA_AND3</type>
<position>-72.5,22.5</position>
<input>
<ID>IN_0</ID>1169 </input>
<input>
<ID>IN_1</ID>1170 </input>
<input>
<ID>IN_2</ID>1171 </input>
<output>
<ID>OUT</ID>1061 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1004</ID>
<type>AA_AND2</type>
<position>-136.5,8</position>
<input>
<ID>IN_0</ID>1152 </input>
<input>
<ID>IN_1</ID>1149 </input>
<output>
<ID>OUT</ID>1141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1009</ID>
<type>DA_FROM</type>
<position>-135.5,0.5</position>
<input>
<ID>IN_0</ID>1146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /T0</lparam></gate>
<gate>
<ID>1016</ID>
<type>DA_FROM</type>
<position>-149.5,3.5</position>
<input>
<ID>IN_0</ID>1150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGI</lparam></gate>
<gate>
<ID>1017</ID>
<type>DA_FROM</type>
<position>-149.5,5.5</position>
<input>
<ID>IN_0</ID>1151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID FGO</lparam></gate>
<gate>
<ID>1018</ID>
<type>DA_FROM</type>
<position>-142.5,9</position>
<input>
<ID>IN_0</ID>1152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IEN</lparam></gate>
<gate>
<ID>1023</ID>
<type>AA_AND3</type>
<position>-72.5,46.5</position>
<input>
<ID>IN_0</ID>1163 </input>
<input>
<ID>IN_1</ID>1164 </input>
<input>
<ID>IN_2</ID>1165 </input>
<output>
<ID>OUT</ID>1155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>1032</ID>
<type>DA_FROM</type>
<position>-78.5,46.5</position>
<input>
<ID>IN_0</ID>1164 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>1033</ID>
<type>DA_FROM</type>
<position>-78.5,44.5</position>
<input>
<ID>IN_0</ID>1165 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Cout</lparam></gate>
<gate>
<ID>1012</ID>
<type>AA_LABEL</type>
<position>-115.5,120.5</position>
<gparam>LABEL_TEXT AC and DR = 0</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1037</ID>
<type>DA_FROM</type>
<position>-78.5,24.5</position>
<input>
<ID>IN_0</ID>1169 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>1038</ID>
<type>DA_FROM</type>
<position>-78.5,22.5</position>
<input>
<ID>IN_0</ID>1170 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T5</lparam></gate>
<gate>
<ID>1039</ID>
<type>DA_FROM</type>
<position>-78.5,20.5</position>
<input>
<ID>IN_0</ID>1171 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /Cout</lparam></gate>
<gate>
<ID>1044</ID>
<type>DA_FROM</type>
<position>-78.5,15.5</position>
<input>
<ID>IN_0</ID>1147 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR10</lparam></gate>
<gate>
<ID>1050</ID>
<type>AA_AND2</type>
<position>80,14.5</position>
<input>
<ID>IN_0</ID>1181 </input>
<input>
<ID>IN_1</ID>1182 </input>
<output>
<ID>OUT</ID>1178 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1052</ID>
<type>DA_FROM</type>
<position>74,15.5</position>
<input>
<ID>IN_0</ID>1181 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1058</ID>
<type>AE_OR2</type>
<position>68,9</position>
<input>
<ID>IN_0</ID>1185 </input>
<input>
<ID>IN_1</ID>1186 </input>
<output>
<ID>OUT</ID>1184 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1063</ID>
<type>DA_FROM</type>
<position>74,11</position>
<input>
<ID>IN_0</ID>1187 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T4</lparam></gate>
<gate>
<ID>70</ID>
<type>DA_FROM</type>
<position>-137,51.5</position>
<input>
<ID>IN_0</ID>80 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>1066</ID>
<type>DA_FROM</type>
<position>74,6.5</position>
<input>
<ID>IN_0</ID>1190 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T6</lparam></gate>
<gate>
<ID>350</ID>
<type>AE_OR3</type>
<position>-29,109.5</position>
<input>
<ID>IN_0</ID>905 </input>
<input>
<ID>IN_1</ID>902 </input>
<input>
<ID>IN_2</ID>24 </input>
<output>
<ID>OUT</ID>906 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>675</ID>
<type>BE_JKFF_LOW</type>
<position>-116.5,18.5</position>
<input>
<ID>J</ID>937 </input>
<input>
<ID>K</ID>940 </input>
<output>
<ID>Q</ID>909 </output>
<input>
<ID>clock</ID>936 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>758</ID>
<type>DE_TO</type>
<position>-110.5,20.5</position>
<input>
<ID>IN_0</ID>909 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID s</lparam></gate>
<gate>
<ID>760</ID>
<type>DA_FROM</type>
<position>-122.5,18.5</position>
<input>
<ID>IN_0</ID>936 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID clk</lparam></gate>
<gate>
<ID>773</ID>
<type>DA_FROM</type>
<position>-122.5,20.5</position>
<input>
<ID>IN_0</ID>937 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>826</ID>
<type>AA_AND2</type>
<position>-123.5,15</position>
<input>
<ID>IN_0</ID>943 </input>
<input>
<ID>IN_1</ID>949 </input>
<output>
<ID>OUT</ID>940 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>889</ID>
<type>DA_FROM</type>
<position>-129.5,14</position>
<input>
<ID>IN_0</ID>949 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR0</lparam></gate>
<gate>
<ID>930</ID>
<type>AE_OR2</type>
<position>31,109</position>
<input>
<ID>IN_0</ID>956 </input>
<input>
<ID>IN_1</ID>955 </input>
<output>
<ID>OUT</ID>954 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>942</ID>
<type>DA_FROM</type>
<position>25,110</position>
<input>
<ID>IN_0</ID>956 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>947</ID>
<type>DA_FROM</type>
<position>66,110</position>
<input>
<ID>IN_0</ID>958 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T1</lparam></gate>
<gate>
<ID>960</ID>
<type>AA_AND2</type>
<position>72,111</position>
<input>
<ID>IN_0</ID>957 </input>
<input>
<ID>IN_1</ID>958 </input>
<output>
<ID>OUT</ID>966 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>966</ID>
<type>AE_OR2</type>
<position>79,114</position>
<input>
<ID>IN_0</ID>1003 </input>
<input>
<ID>IN_1</ID>966 </input>
<output>
<ID>OUT</ID>1035 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>618</ID>
<type>DA_FROM</type>
<position>127,19</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID p</lparam></gate>
<gate>
<ID>977</ID>
<type>DA_FROM</type>
<position>73,115</position>
<input>
<ID>IN_0</ID>1003 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID START</lparam></gate>
<gate>
<ID>993</ID>
<type>AA_LABEL</type>
<position>-94.5,67.5</position>
<gparam>LABEL_TEXT Flags & Flip Flops</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1001</ID>
<type>AA_LABEL</type>
<position>-19,36</position>
<gparam>LABEL_TEXT Sequence Counter</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1005</ID>
<type>AA_LABEL</type>
<position>-20,61.5</position>
<gparam>LABEL_TEXT IR Decoder</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1010</ID>
<type>AA_LABEL</type>
<position>14.5,17</position>
<gparam>LABEL_TEXT p and r bits</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1014</ID>
<type>AA_LABEL</type>
<position>-66.5,123</position>
<gparam>LABEL_TEXT ALU Control Signals</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1021</ID>
<type>AA_LABEL</type>
<position>-22,129.5</position>
<gparam>LABEL_TEXT AC Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1045</ID>
<type>AA_LABEL</type>
<position>27.5,77.5</position>
<gparam>LABEL_TEXT Memory Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1053</ID>
<type>AA_LABEL</type>
<position>79.5,133.5</position>
<gparam>LABEL_TEXT PC Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1062</ID>
<type>AA_LABEL</type>
<position>132.5,81.5</position>
<gparam>LABEL_TEXT IR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>1068</ID>
<type>AA_LABEL</type>
<position>133.5,58.5</position>
<gparam>LABEL_TEXT TR Control</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>775</ID>
<type>AA_AND2</type>
<position>-83,5.5</position>
<input>
<ID>IN_0</ID>1158 </input>
<input>
<ID>IN_1</ID>1160 </input>
<output>
<ID>OUT</ID>1154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>811</ID>
<type>AA_AND2</type>
<position>-83,0.5</position>
<input>
<ID>IN_0</ID>1159 </input>
<input>
<ID>IN_1</ID>1172 </input>
<output>
<ID>OUT</ID>1157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>834</ID>
<type>DA_FROM</type>
<position>-89,6.5</position>
<input>
<ID>IN_0</ID>1158 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR7</lparam></gate>
<gate>
<ID>990</ID>
<type>DA_FROM</type>
<position>-94,4.5</position>
<input>
<ID>IN_0</ID>1161 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo0</lparam></gate>
<gate>
<ID>1006</ID>
<type>DA_FROM</type>
<position>-89,37.5</position>
<input>
<ID>IN_0</ID>1176 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID /E</lparam></gate>
<gate>
<ID>1011</ID>
<type>DA_FROM</type>
<position>-89,29.5</position>
<input>
<ID>IN_0</ID>1196 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID IR6</lparam></gate>
<gate>
<ID>1022</ID>
<type>DA_FROM</type>
<position>-89,27.5</position>
<input>
<ID>IN_0</ID>1202 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID ACo15</lparam></gate>
<gate>
<ID>1028</ID>
<type>AA_AND2</type>
<position>-83,33.5</position>
<input>
<ID>IN_0</ID>1195 </input>
<input>
<ID>IN_1</ID>1203 </input>
<output>
<ID>OUT</ID>1193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>5</ID>
<type>AE_OR2</type>
<position>-123.5,54</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>90</ID>
<type>DA_FROM</type>
<position>-137,49.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>-129.5,-2</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID R</lparam></gate>
<gate>
<ID>106</ID>
<type>DA_FROM</type>
<position>-129.5,-4</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID T2</lparam></gate>
<wire>
<ID>1103 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,66,35,66</points>
<connection>
<GID>941</GID>
<name>OUT</name></connection>
<connection>
<GID>768</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1039 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>74.5,69.5,75.5,69.5</points>
<connection>
<GID>921</GID>
<name>IN_0</name></connection>
<connection>
<GID>901</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,19,-26,19</points>
<connection>
<GID>138</GID>
<name>IN_3</name></connection>
<connection>
<GID>7</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>950 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,84.5,-115,84.5</points>
<connection>
<GID>849</GID>
<name>IN_0</name></connection>
<connection>
<GID>807</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>713 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>-120.5,31.5,-119.5,31.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<connection>
<GID>319</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1043 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>74.5,78.5,75.5,78.5</points>
<connection>
<GID>917</GID>
<name>IN_0</name></connection>
<connection>
<GID>900</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>408 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,24,-17,24</points>
<connection>
<GID>138</GID>
<name>OUT_8</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>609 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,51,-18,51</points>
<connection>
<GID>46</GID>
<name>OUT_4</name></connection>
<connection>
<GID>160</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1078 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,118,-25,118</points>
<connection>
<GID>833</GID>
<name>IN_0</name></connection>
<connection>
<GID>777</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>959 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,117,-63,117</points>
<connection>
<GID>748</GID>
<name>IN_0</name></connection>
<connection>
<GID>836</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>911 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,104,-108,107</points>
<connection>
<GID>774</GID>
<name>OUT</name></connection>
<intersection>107 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,107,-107,107</points>
<connection>
<GID>776</GID>
<name>IN_1</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>1030 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,99.5,75.5,99.5</points>
<connection>
<GID>896</GID>
<name>IN_0</name></connection>
<connection>
<GID>908</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>337 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71,85,-70,85</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<connection>
<GID>281</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>636 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,52,-12.5,52</points>
<connection>
<GID>46</GID>
<name>OUT_5</name></connection>
<connection>
<GID>168</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>923 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,50,21,50</points>
<connection>
<GID>792</GID>
<name>IN_1</name></connection>
<connection>
<GID>779</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>406 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,18,-17,18</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_2</name></connection>
<intersection>-18.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-18.5,9,-18.5,18</points>
<intersection>9 15</intersection>
<intersection>18 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-18.5,9,-18,9</points>
<connection>
<GID>997</GID>
<name>IN_0</name></connection>
<intersection>-18.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>683 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,54,-12.5,54</points>
<connection>
<GID>46</GID>
<name>OUT_7</name></connection>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-18.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-18.5,54,-18.5,56.5</points>
<intersection>54 1</intersection>
<intersection>56.5 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-18.5,56.5,-17.5,56.5</points>
<connection>
<GID>783</GID>
<name>IN_0</name></connection>
<intersection>-18.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>319 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-31,22,-31,24</points>
<connection>
<GID>7</GID>
<name>count_enable</name></connection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33,24,-31,24</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>-31 0</intersection></hsegment></shape></wire>
<wire>
<ID>1196 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,29.5,-86,29.5</points>
<connection>
<GID>1029</GID>
<name>IN_0</name></connection>
<connection>
<GID>1011</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,10,13,10</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-135,51.5,-134,51.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1132 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,59.5,-75,62</points>
<connection>
<GID>986</GID>
<name>IN_0</name></connection>
<intersection>62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76,62,-73,62</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<connection>
<GID>982</GID>
<name>IN_0</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>322 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,95,-63,95</points>
<connection>
<GID>259</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1113 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,58.5,21,58.5</points>
<connection>
<GID>958</GID>
<name>IN_0</name></connection>
<connection>
<GID>946</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>964 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,111.5,-63,111.5</points>
<connection>
<GID>750</GID>
<name>IN_0</name></connection>
<connection>
<GID>841</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>999 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,106,-63,106</points>
<connection>
<GID>752</GID>
<name>IN_0</name></connection>
<connection>
<GID>871</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1054 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,58.5,62,58.5</points>
<connection>
<GID>933</GID>
<name>IN_0</name></connection>
<connection>
<GID>935</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,22,-17,22</points>
<connection>
<GID>138</GID>
<name>OUT_6</name></connection>
<connection>
<GID>228</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-135,49.5,-134,49.5</points>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<connection>
<GID>90</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>12,12,13,12</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1074 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,120,-25.5,122.5</points>
<intersection>120 3</intersection>
<intersection>122.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-26,122.5,-25.5,122.5</points>
<connection>
<GID>814</GID>
<name>OUT</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-25.5,120,-25,120</points>
<connection>
<GID>777</GID>
<name>IN_0</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-127,50.5,-127,53</points>
<intersection>50.5 2</intersection>
<intersection>53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-127,53,-126.5,53</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>-127 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-128,50.5,-127,50.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<intersection>-127 0</intersection></hsegment></shape></wire>
<wire>
<ID>896 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>67.5,125.5,68.5,125.5</points>
<connection>
<GID>751</GID>
<name>IN_0</name></connection>
<connection>
<GID>741</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,19,-10.5,19</points>
<connection>
<GID>138</GID>
<name>OUT_3</name></connection>
<connection>
<GID>175</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>499 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,49,-26.5,50</points>
<intersection>49 1</intersection>
<intersection>50 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26.5,49,-26,49</points>
<connection>
<GID>46</GID>
<name>IN_2</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-27.5,50,-26.5,50</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,2,13,2</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1173 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,40.5,-75.5,40.5</points>
<connection>
<GID>994</GID>
<name>IN_0</name></connection>
<connection>
<GID>1026</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>904 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,12.5,-75.5,12.5</points>
<connection>
<GID>1040</GID>
<name>IN_0</name></connection>
<connection>
<GID>377</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1120 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,39.5,-126.5,39.5</points>
<connection>
<GID>965</GID>
<name>IN_1</name></connection>
<connection>
<GID>968</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>941 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,38.5,27.5,42</points>
<intersection>38.5 9</intersection>
<intersection>42 10</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>27,38.5,27.5,38.5</points>
<connection>
<GID>809</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>27.5,42,28,42</points>
<connection>
<GID>815</GID>
<name>IN_2</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>411 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,16,-17,16</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-19.5 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-19.5,13,-19.5,16</points>
<intersection>13 15</intersection>
<intersection>16 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-19.5,13,-15,13</points>
<connection>
<GID>995</GID>
<name>IN_0</name></connection>
<intersection>-19.5 14</intersection></hsegment></shape></wire>
<wire>
<ID>917 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,105.5,-115,105.5</points>
<connection>
<GID>774</GID>
<name>IN_2</name></connection>
<connection>
<GID>793</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1096 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,36.5,13,36.5</points>
<connection>
<GID>812</GID>
<name>IN_0</name></connection>
<connection>
<GID>925</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1097 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,34.5,13,34.5</points>
<connection>
<GID>813</GID>
<name>IN_0</name></connection>
<connection>
<GID>925</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>891 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,86.5,21,86.5</points>
<connection>
<GID>739</GID>
<name>IN_0</name></connection>
<connection>
<GID>649</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1098 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,32.5,13,32.5</points>
<connection>
<GID>926</GID>
<name>IN_0</name></connection>
<connection>
<GID>925</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,18,-26,18</points>
<connection>
<GID>138</GID>
<name>IN_2</name></connection>
<connection>
<GID>7</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>922 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,48,21,48</points>
<connection>
<GID>792</GID>
<name>IN_2</name></connection>
<connection>
<GID>785</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1099 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,30.5,13,30.5</points>
<connection>
<GID>928</GID>
<name>IN_0</name></connection>
<connection>
<GID>925</GID>
<name>IN_3</name></connection></hsegment></shape></wire>
<wire>
<ID>1095 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,33.5,20.5,37.5</points>
<intersection>33.5 2</intersection>
<intersection>37.5 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>20,33.5,20.5,33.5</points>
<connection>
<GID>925</GID>
<name>OUT</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>20.5,37.5,21,37.5</points>
<connection>
<GID>809</GID>
<name>IN_1</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1046 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,62.5,75.5,62.5</points>
<connection>
<GID>902</GID>
<name>IN_2</name></connection>
<connection>
<GID>923</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>688 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>-120.5,44,-119.5,44</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<connection>
<GID>311</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,27,-10.5,27</points>
<connection>
<GID>138</GID>
<name>OUT_11</name></connection>
<connection>
<GID>236</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1006 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,89.5,-115,89.5</points>
<connection>
<GID>837</GID>
<name>IN_0</name></connection>
<connection>
<GID>805</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,31,-10.5,31</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_15</name></connection></hsegment></shape></wire>
<wire>
<ID>942 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,50,27.5,50</points>
<connection>
<GID>792</GID>
<name>OUT</name></connection>
<intersection>27.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>27.5,46,27.5,50</points>
<intersection>46 11</intersection>
<intersection>50 1</intersection></vsegment>
<hsegment>
<ID>11</ID>
<points>27.5,46,28,46</points>
<connection>
<GID>815</GID>
<name>IN_0</name></connection>
<intersection>27.5 10</intersection></hsegment></shape></wire>
<wire>
<ID>1143 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,17.5,-75.5,17.5</points>
<connection>
<GID>759</GID>
<name>IN_0</name></connection>
<connection>
<GID>757</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>324 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,88.5,-70,88.5</points>
<connection>
<GID>275</GID>
<name>IN_0</name></connection>
<connection>
<GID>273</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,39.5,-86,39.5</points>
<connection>
<GID>1003</GID>
<name>IN_0</name></connection>
<connection>
<GID>1024</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>910 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,109,-108,112</points>
<connection>
<GID>770</GID>
<name>OUT</name></connection>
<intersection>109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,109,-107,109</points>
<connection>
<GID>776</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>412 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,30,-17,30</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_14</name></connection></hsegment></shape></wire>
<wire>
<ID>934 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101,108,-100,108</points>
<connection>
<GID>776</GID>
<name>OUT</name></connection>
<connection>
<GID>803</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1102 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,45,21,45</points>
<connection>
<GID>939</GID>
<name>IN_0</name></connection>
<connection>
<GID>932</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>409 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,20,-17,20</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_4</name></connection></hsegment></shape></wire>
<wire>
<ID>791 </ID>
<shape>
<hsegment>
<ID>13</ID>
<points>20,105,21,105</points>
<connection>
<GID>548</GID>
<name>IN_1</name></connection>
<connection>
<GID>574</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>242 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-30,9.5,-30,13</points>
<connection>
<GID>7</GID>
<name>clear</name></connection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,9.5,-30,9.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>-30 0</intersection></hsegment></shape></wire>
<wire>
<ID>1201 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,28.5,-69,37.5</points>
<intersection>28.5 1</intersection>
<intersection>37.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,28.5,-68,28.5</points>
<connection>
<GID>1020</GID>
<name>IN_1</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,37.5,-69,37.5</points>
<connection>
<GID>1026</GID>
<name>OUT</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>205 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,11.5,-32,13</points>
<connection>
<GID>7</GID>
<name>clock</name></connection>
<intersection>11.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-33.5,11.5,-32,11.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>-32 0</intersection></hsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,23,-10.5,23</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_7</name></connection></hsegment></shape></wire>
<wire>
<ID>1073 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,115,-18.5,119</points>
<intersection>115 1</intersection>
<intersection>119 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-18.5,115,-18,115</points>
<connection>
<GID>549</GID>
<name>IN_0</name></connection>
<intersection>-18.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19,119,-18.5,119</points>
<connection>
<GID>777</GID>
<name>OUT</name></connection>
<intersection>-18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>924 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,114.5,-115,114.5</points>
<connection>
<GID>770</GID>
<name>IN_1</name></connection>
<connection>
<GID>780</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,16,-26,16</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1021 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,71.5,89.5,80.5</points>
<intersection>71.5 1</intersection>
<intersection>80.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,71.5,89.5,71.5</points>
<connection>
<GID>901</GID>
<name>OUT</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,80.5,97.5,80.5</points>
<connection>
<GID>880</GID>
<name>IN_6</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>534 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26.5,46,-26.5,47</points>
<intersection>46 1</intersection>
<intersection>47 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-27.5,46,-26.5,46</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26.5,47,-26,47</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>-26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,17,-26,17</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,44,28,44</points>
<connection>
<GID>932</GID>
<name>OUT</name></connection>
<connection>
<GID>815</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>939 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,44,35,44</points>
<connection>
<GID>769</GID>
<name>IN_0</name></connection>
<connection>
<GID>815</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1044 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,114,-25,114</points>
<connection>
<GID>623</GID>
<name>IN_0</name></connection>
<connection>
<GID>696</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,17,-10.5,17</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_1</name></connection>
<intersection>-19 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>-19,11,-19,17</points>
<intersection>11 15</intersection>
<intersection>17 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-19,11,-16.5,11</points>
<connection>
<GID>996</GID>
<name>IN_0</name></connection>
<intersection>-19 14</intersection></hsegment></shape></wire>
<wire>
<ID>1092 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>127.5,48,128.5,48</points>
<connection>
<GID>895</GID>
<name>IN_0</name></connection>
<connection>
<GID>897</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>407 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,26,-17,26</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_10</name></connection></hsegment></shape></wire>
<wire>
<ID>410 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,28,-17,28</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_12</name></connection></hsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,29,-10.5,29</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_13</name></connection></hsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,21,-10.5,21</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1187 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,11,77,11</points>
<connection>
<GID>1056</GID>
<name>IN_0</name></connection>
<connection>
<GID>1063</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1010 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,9.5,-86,9.5</points>
<connection>
<GID>1042</GID>
<name>IN_0</name></connection>
<connection>
<GID>671</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>23 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-67,57.5,-66,57.5</points>
<connection>
<GID>317</GID>
<name>IN_0</name></connection>
<connection>
<GID>158</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,25,-10.5,25</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>OUT_9</name></connection></hsegment></shape></wire>
<wire>
<ID>1086 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,78,-19,78</points>
<connection>
<GID>888</GID>
<name>IN_0</name></connection>
<connection>
<GID>887</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>967 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,94.5,-115,94.5</points>
<connection>
<GID>823</GID>
<name>IN_0</name></connection>
<connection>
<GID>805</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,32.5,-86,32.5</points>
<connection>
<GID>1034</GID>
<name>IN_0</name></connection>
<connection>
<GID>1028</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>898 </ID>
<shape>
<hsegment>
<ID>18</ID>
<points>120,102,121,102</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>962 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,112.5,-70,112.5</points>
<connection>
<GID>841</GID>
<name>IN_0</name></connection>
<connection>
<GID>842</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>963 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,110.5,-70,110.5</points>
<connection>
<GID>841</GID>
<name>IN_1</name></connection>
<connection>
<GID>843</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1174 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,38.5,-75.5,38.5</points>
<connection>
<GID>1026</GID>
<name>IN_1</name></connection>
<connection>
<GID>1024</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>350 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,84,-63,84</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<connection>
<GID>281</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1193 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,33.5,-78,36.5</points>
<intersection>33.5 2</intersection>
<intersection>36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,36.5,-75.5,36.5</points>
<connection>
<GID>1026</GID>
<name>IN_2</name></connection>
<intersection>-78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80,33.5,-78,33.5</points>
<connection>
<GID>1028</GID>
<name>OUT</name></connection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>1194 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,28.5,-77.5,34.5</points>
<intersection>28.5 2</intersection>
<intersection>34.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,34.5,-75.5,34.5</points>
<connection>
<GID>1026</GID>
<name>IN_3</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80,28.5,-77.5,28.5</points>
<connection>
<GID>1029</GID>
<name>OUT</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1130 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,59.5,-66.5,61</points>
<intersection>59.5 1</intersection>
<intersection>61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-66.5,59.5,-66,59.5</points>
<connection>
<GID>158</GID>
<name>J</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-67,61,-66.5,61</points>
<connection>
<GID>982</GID>
<name>OUT</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>954 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,109,35,109</points>
<connection>
<GID>930</GID>
<name>OUT</name></connection>
<connection>
<GID>592</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1131 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-66.5,54,-66.5,55.5</points>
<intersection>54 1</intersection>
<intersection>55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-67,54,-66.5,54</points>
<connection>
<GID>984</GID>
<name>OUT</name></connection>
<intersection>-66.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-66.5,55.5,-66,55.5</points>
<connection>
<GID>158</GID>
<name>K</name></connection>
<intersection>-66.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>733 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,59.5,-111.5,59.5</points>
<connection>
<GID>302</GID>
<name>Q</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection>
<intersection>-112.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-112.5,59.5,-112.5,61</points>
<connection>
<GID>308</GID>
<name>N_in2</name></connection>
<intersection>59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>886 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-60,59.5,-58,59.5</points>
<connection>
<GID>158</GID>
<name>Q</name></connection>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>-59 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-59,59.5,-59,61</points>
<connection>
<GID>847</GID>
<name>N_in2</name></connection>
<intersection>59.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-60,55.5,-58,55.5</points>
<connection>
<GID>158</GID>
<name>nQ</name></connection>
<connection>
<GID>68</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1180 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,20,77,20</points>
<connection>
<GID>819</GID>
<name>IN_0</name></connection>
<connection>
<GID>875</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,8,13,8</points>
<connection>
<GID>51</GID>
<name>IN_2</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1002 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,23,64,23</points>
<connection>
<GID>821</GID>
<name>IN_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,18,77,18</points>
<connection>
<GID>819</GID>
<name>IN_1</name></connection>
<connection>
<GID>820</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>948 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,19,84,19</points>
<connection>
<GID>819</GID>
<name>OUT</name></connection>
<intersection>84 14</intersection></hsegment>
<vsegment>
<ID>14</ID>
<points>84,8.5,84,19</points>
<intersection>8.5 15</intersection>
<intersection>19 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>84,8.5,84.5,8.5</points>
<connection>
<GID>824</GID>
<name>IN_0</name></connection>
<intersection>84 14</intersection></hsegment></shape></wire>
<wire>
<ID>1115 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,33.5,-119.5,33.5</points>
<connection>
<GID>319</GID>
<name>J</name></connection>
<connection>
<GID>961</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>938 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,11.5,-86,11.5</points>
<connection>
<GID>1041</GID>
<name>IN_0</name></connection>
<connection>
<GID>671</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>978 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,83.5,-115,83.5</points>
<connection>
<GID>807</GID>
<name>IN_6</name></connection>
<connection>
<GID>850</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1155 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,30.5,-68.5,46.5</points>
<intersection>30.5 1</intersection>
<intersection>46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,30.5,-68,30.5</points>
<connection>
<GID>1020</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,46.5,-68.5,46.5</points>
<connection>
<GID>1023</GID>
<name>OUT</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1153 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,28,-61.5,29.5</points>
<intersection>28 1</intersection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61.5,28,-61,28</points>
<connection>
<GID>297</GID>
<name>J</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62,29.5,-61.5,29.5</points>
<connection>
<GID>1020</GID>
<name>OUT</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1101 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,43,21,43</points>
<connection>
<GID>932</GID>
<name>IN_1</name></connection>
<connection>
<GID>771</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>500 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27.5,48,-26,48</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>610 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,47,-18,47</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>661 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,48,-12.5,48</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_1</name></connection></hsegment></shape></wire>
<wire>
<ID>635 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,49,-18,49</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_2</name></connection></hsegment></shape></wire>
<wire>
<ID>682 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,50,-12.5,50</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_3</name></connection></hsegment></shape></wire>
<wire>
<ID>535 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,53,-18,53</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>46</GID>
<name>OUT_6</name></connection></hsegment></shape></wire>
<wire>
<ID>1159 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,1.5,-86,1.5</points>
<connection>
<GID>877</GID>
<name>IN_0</name></connection>
<connection>
<GID>811</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1005 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,91.5,-115,91.5</points>
<connection>
<GID>805</GID>
<name>IN_6</name></connection>
<connection>
<GID>828</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1184 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71,9,77,9</points>
<connection>
<GID>1056</GID>
<name>IN_1</name></connection>
<connection>
<GID>1058</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1183 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,6.5,83,10</points>
<connection>
<GID>1056</GID>
<name>OUT</name></connection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,6.5,84.5,6.5</points>
<connection>
<GID>824</GID>
<name>IN_2</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>349 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,83,-70,83</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<connection>
<GID>281</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1035 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>82,114,83,114</points>
<connection>
<GID>646</GID>
<name>IN_0</name></connection>
<connection>
<GID>966</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1135 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-84,58.5,-83,58.5</points>
<connection>
<GID>988</GID>
<name>IN_0</name></connection>
<connection>
<GID>980</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1036 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,85.5,75.5,85.5</points>
<connection>
<GID>899</GID>
<name>IN_1</name></connection>
<connection>
<GID>914</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,-0.5,-111.5,-0.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<connection>
<GID>289</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>1089 </ID>
<shape>
<hsegment>
<ID>9</ID>
<points>127.5,54,128.5,54</points>
<connection>
<GID>891</GID>
<name>IN_0</name></connection>
<connection>
<GID>892</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1091 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>134.5,53,135.5,53</points>
<connection>
<GID>892</GID>
<name>OUT</name></connection>
<connection>
<GID>764</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>914 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13.5,56.5,-12.5,56.5</points>
<connection>
<GID>781</GID>
<name>IN_0</name></connection>
<connection>
<GID>783</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>929 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,106.5,-115,106.5</points>
<connection>
<GID>791</GID>
<name>IN_0</name></connection>
<connection>
<GID>774</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1053 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,56.5,62,56.5</points>
<connection>
<GID>933</GID>
<name>IN_1</name></connection>
<connection>
<GID>936</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>714 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,33.5,-111.5,33.5</points>
<connection>
<GID>319</GID>
<name>Q</name></connection>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>-112.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-112.5,33.5,-112.5,35</points>
<connection>
<GID>349</GID>
<name>N_in2</name></connection>
<intersection>33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>1052 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,56,68,57.5</points>
<connection>
<GID>933</GID>
<name>OUT</name></connection>
<intersection>56 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68,56,68.5,56</points>
<connection>
<GID>931</GID>
<name>IN_0</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>1163 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-76.5,48.5,-75.5,48.5</points>
<connection>
<GID>1031</GID>
<name>IN_0</name></connection>
<connection>
<GID>1023</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1127 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-120,59.5,-120,61</points>
<intersection>59.5 1</intersection>
<intersection>61 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-120,59.5,-119.5,59.5</points>
<connection>
<GID>302</GID>
<name>J</name></connection>
<intersection>-120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-120.5,61,-120,61</points>
<connection>
<GID>975</GID>
<name>OUT</name></connection>
<intersection>-120 0</intersection></hsegment></shape></wire>
<wire>
<ID>1087 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,77,-12,77</points>
<connection>
<GID>731</GID>
<name>IN_0</name></connection>
<connection>
<GID>888</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-120,54,-120,55.5</points>
<intersection>54 2</intersection>
<intersection>55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-120,55.5,-119.5,55.5</points>
<connection>
<GID>302</GID>
<name>K</name></connection>
<intersection>-120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-120.5,54,-120,54</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-120 0</intersection></hsegment></shape></wire>
<wire>
<ID>470 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,57.5,-119.5,57.5</points>
<connection>
<GID>302</GID>
<name>clock</name></connection>
<connection>
<GID>301</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>469 </ID>
<shape>
<hsegment>
<ID>3</ID>
<points>-113.5,55.5,-111.5,55.5</points>
<connection>
<GID>302</GID>
<name>nQ</name></connection>
<connection>
<GID>309</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1138 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12.5,11,-11.5,11</points>
<connection>
<GID>999</GID>
<name>IN_0</name></connection>
<connection>
<GID>996</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>443 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-62,26,-61,26</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>1139 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14,9,-13,9</points>
<connection>
<GID>997</GID>
<name>OUT_0</name></connection>
<connection>
<GID>1000</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,99.5,-70,99.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<hsegment>
<ID>7</ID>
<points>-120.5,1.5,-119.5,1.5</points>
<connection>
<GID>289</GID>
<name>clock</name></connection>
<connection>
<GID>287</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1058 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,34,135.5,34</points>
<connection>
<GID>762</GID>
<name>IN_0</name></connection>
<connection>
<GID>983</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>734 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,128.5,20.5,128.5</points>
<connection>
<GID>403</GID>
<name>OUT</name></connection>
<intersection>20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>20.5,127,20.5,128.5</points>
<intersection>127 4</intersection>
<intersection>128.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>20.5,127,21,127</points>
<connection>
<GID>376</GID>
<name>IN_0</name></connection>
<intersection>20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>740 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,125,21,125</points>
<connection>
<GID>457</GID>
<name>IN_0</name></connection>
<connection>
<GID>376</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>739 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,125,27.5,126</points>
<intersection>125 1</intersection>
<intersection>126 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,125,28,125</points>
<connection>
<GID>430</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,126,27.5,126</points>
<connection>
<GID>376</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>882 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,100,35,100</points>
<connection>
<GID>595</GID>
<name>OUT</name></connection>
<connection>
<GID>553</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>880 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,101,28,101</points>
<connection>
<GID>617</GID>
<name>IN_0</name></connection>
<connection>
<GID>595</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>735 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,124,35,124</points>
<connection>
<GID>430</GID>
<name>OUT</name></connection>
<connection>
<GID>577</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71,96,-70,96</points>
<connection>
<GID>261</GID>
<name>IN_0</name></connection>
<connection>
<GID>263</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1090 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,52,128.5,52</points>
<connection>
<GID>892</GID>
<name>IN_1</name></connection>
<connection>
<GID>893</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>883 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,89.5,35,89.5</points>
<connection>
<GID>619</GID>
<name>OUT</name></connection>
<connection>
<GID>596</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1008 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104.5,82,105.5,82</points>
<connection>
<GID>622</GID>
<name>IN_0</name></connection>
<connection>
<GID>880</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1161 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92,4.5,-91,4.5</points>
<connection>
<GID>981</GID>
<name>IN_0</name></connection>
<connection>
<GID>990</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>981 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,87.5,-115,87.5</points>
<connection>
<GID>807</GID>
<name>IN_1</name></connection>
<connection>
<GID>844</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1160 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,4.5,-86,4.5</points>
<connection>
<GID>981</GID>
<name>OUT_0</name></connection>
<connection>
<GID>775</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1049 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,83.5,70.5,83.5</points>
<connection>
<GID>927</GID>
<name>IN_0</name></connection>
<connection>
<GID>929</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>900 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,126.5,82.5,126.5</points>
<connection>
<GID>644</GID>
<name>IN_0</name></connection>
<connection>
<GID>743</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1037 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,71.5,75.5,71.5</points>
<connection>
<GID>901</GID>
<name>IN_1</name></connection>
<connection>
<GID>915</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>687 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,42,-111.5,42</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<connection>
<GID>311</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>890 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,88.5,21,88.5</points>
<connection>
<GID>723</GID>
<name>IN_0</name></connection>
<connection>
<GID>649</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1067 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>81.5,44.5,82.5,44.5</points>
<connection>
<GID>650</GID>
<name>IN_0</name></connection>
<connection>
<GID>952</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>707 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,46,-111.5,46</points>
<connection>
<GID>311</GID>
<name>Q</name></connection>
<connection>
<GID>313</GID>
<name>IN_0</name></connection>
<intersection>-112.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-112.5,46,-112.5,47.5</points>
<connection>
<GID>314</GID>
<name>N_in2</name></connection>
<intersection>46 1</intersection></vsegment></shape></wire>
<wire>
<ID>21 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,110.5,135.5,110.5</points>
<connection>
<GID>698</GID>
<name>IN_0</name></connection>
<connection>
<GID>50</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1107 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,62.5,20.5,62.5</points>
<connection>
<GID>951</GID>
<name>OUT</name></connection>
<intersection>20.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>20.5,62.5,20.5,65</points>
<intersection>62.5 1</intersection>
<intersection>65 8</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>20.5,65,21,65</points>
<connection>
<GID>943</GID>
<name>IN_1</name></connection>
<intersection>20.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>930 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,128,135.5,128</points>
<connection>
<GID>701</GID>
<name>IN_0</name></connection>
<connection>
<GID>800</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1009 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134,99,135.5,99</points>
<connection>
<GID>722</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,10,65,10</points>
<connection>
<GID>1060</GID>
<name>IN_0</name></connection>
<connection>
<GID>1058</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>85 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>136,18,137,18</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>932 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,102.5,-115,102.5</points>
<connection>
<GID>774</GID>
<name>IN_6</name></connection>
<connection>
<GID>797</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1081 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,85,-12,85</points>
<connection>
<GID>727</GID>
<name>IN_0</name></connection>
<connection>
<GID>1075</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1176 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,37.5,-86,37.5</points>
<connection>
<GID>1024</GID>
<name>IN_1</name></connection>
<connection>
<GID>1006</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>997 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71,107,-70,107</points>
<connection>
<GID>872</GID>
<name>IN_0</name></connection>
<connection>
<GID>871</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>885 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,87.5,27.5,88.5</points>
<intersection>87.5 2</intersection>
<intersection>88.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,88.5,28,88.5</points>
<connection>
<GID>619</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,87.5,27.5,87.5</points>
<connection>
<GID>649</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1064 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,91,-12,91</points>
<connection>
<GID>728</GID>
<name>IN_0</name></connection>
<connection>
<GID>879</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1017 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,113,-11,113</points>
<connection>
<GID>729</GID>
<name>IN_0</name></connection>
<connection>
<GID>549</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1079 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,90,-19,90</points>
<connection>
<GID>882</GID>
<name>IN_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1186 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>64,8,65,8</points>
<connection>
<GID>1059</GID>
<name>IN_0</name></connection>
<connection>
<GID>1058</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1026 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,85.5,90.5,103.5</points>
<intersection>85.5 2</intersection>
<intersection>103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,103.5,90.5,103.5</points>
<connection>
<GID>894</GID>
<name>OUT</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,85.5,97.5,85.5</points>
<connection>
<GID>880</GID>
<name>IN_0</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1004 </ID>
<shape>
<hsegment>
<ID>17</ID>
<points>63,17,64,17</points>
<connection>
<GID>875</GID>
<name>IN_3</name></connection>
<connection>
<GID>876</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1025 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,84.5,90,98.5</points>
<intersection>84.5 2</intersection>
<intersection>98.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,98.5,90,98.5</points>
<connection>
<GID>896</GID>
<name>OUT</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90,84.5,97.5,84.5</points>
<connection>
<GID>880</GID>
<name>IN_1</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>1024 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,83.5,89.5,92.5</points>
<intersection>83.5 2</intersection>
<intersection>92.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,92.5,89.5,92.5</points>
<connection>
<GID>898</GID>
<name>OUT</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89.5,83.5,97.5,83.5</points>
<connection>
<GID>880</GID>
<name>IN_2</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1023 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,82.5,89,85.5</points>
<intersection>82.5 2</intersection>
<intersection>85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,85.5,89,85.5</points>
<connection>
<GID>899</GID>
<name>OUT</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>89,82.5,97.5,82.5</points>
<connection>
<GID>880</GID>
<name>IN_3</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>1019 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,58.5,90.5,78.5</points>
<intersection>58.5 1</intersection>
<intersection>78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,58.5,90.5,58.5</points>
<connection>
<GID>904</GID>
<name>OUT</name></connection>
<intersection>90.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>90.5,78.5,97.5,78.5</points>
<connection>
<GID>880</GID>
<name>IN_4</name></connection>
<intersection>90.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1041 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,80.5,75.5,80.5</points>
<connection>
<GID>900</GID>
<name>IN_0</name></connection>
<connection>
<GID>916</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1020 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,64.5,90,79.5</points>
<intersection>64.5 2</intersection>
<intersection>79.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>90,79.5,97.5,79.5</points>
<connection>
<GID>880</GID>
<name>IN_5</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,64.5,90,64.5</points>
<connection>
<GID>902</GID>
<name>OUT</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>19 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12,0,13,0</points>
<connection>
<GID>65</GID>
<name>IN_2</name></connection>
<connection>
<GID>66</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1022 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89,78.5,89,81.5</points>
<intersection>78.5 2</intersection>
<intersection>81.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>89,81.5,97.5,81.5</points>
<connection>
<GID>880</GID>
<name>IN_7</name></connection>
<intersection>89 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,78.5,89,78.5</points>
<connection>
<GID>900</GID>
<name>OUT</name></connection>
<intersection>89 0</intersection></hsegment></shape></wire>
<wire>
<ID>1192 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83,-1.5,83,3.5</points>
<intersection>-1.5 2</intersection>
<intersection>3.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83,3.5,84.5,3.5</points>
<connection>
<GID>824</GID>
<name>IN_6</name></connection>
<intersection>83 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-1.5,83,-1.5</points>
<connection>
<GID>1070</GID>
<name>IN_0</name></connection>
<intersection>83 0</intersection></hsegment></shape></wire>
<wire>
<ID>1013 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,74.5,135.5,74.5</points>
<connection>
<GID>735</GID>
<name>IN_0</name></connection>
<connection>
<GID>404</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1016 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,69,135.5,69</points>
<connection>
<GID>737</GID>
<name>IN_0</name></connection>
<connection>
<GID>485</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>909 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-113.5,20.5,-112.5,20.5</points>
<connection>
<GID>675</GID>
<name>Q</name></connection>
<connection>
<GID>758</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1088 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>134,40.5,134,41.5</points>
<connection>
<GID>890</GID>
<name>OUT_0</name></connection>
<intersection>41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>134,41.5,135.5,41.5</points>
<connection>
<GID>763</GID>
<name>IN_0</name></connection>
<intersection>134 0</intersection></hsegment></shape></wire>
<wire>
<ID>1189 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,4.5,77,4.5</points>
<connection>
<GID>1067</GID>
<name>IN_0</name></connection>
<connection>
<GID>1065</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>980 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,85.5,-115,85.5</points>
<connection>
<GID>807</GID>
<name>IN_3</name></connection>
<connection>
<GID>848</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1129 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,86,-19,86</points>
<connection>
<GID>1075</GID>
<name>IN_0</name></connection>
<connection>
<GID>987</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1084 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,82,-19.5,84</points>
<intersection>82 2</intersection>
<intersection>84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19.5,84,-19,84</points>
<connection>
<GID>1075</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-20,82,-19.5,82</points>
<connection>
<GID>885</GID>
<name>OUT</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>912 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,115.5,-115,115.5</points>
<connection>
<GID>770</GID>
<name>IN_0</name></connection>
<connection>
<GID>778</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1065 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,41.5,69,41.5</points>
<connection>
<GID>944</GID>
<name>IN_1</name></connection>
<connection>
<GID>950</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>916 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,113.5,-115,113.5</points>
<connection>
<GID>770</GID>
<name>IN_2</name></connection>
<connection>
<GID>782</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>926 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,112.5,-115,112.5</points>
<connection>
<GID>770</GID>
<name>IN_3</name></connection>
<connection>
<GID>784</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>921 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,108.5,-115,108.5</points>
<connection>
<GID>770</GID>
<name>IN_4</name></connection>
<connection>
<GID>789</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>915 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,109.5,-115,109.5</points>
<connection>
<GID>770</GID>
<name>IN_5</name></connection>
<connection>
<GID>788</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>927 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,110.5,-115,110.5</points>
<connection>
<GID>770</GID>
<name>IN_6</name></connection>
<connection>
<GID>787</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>913 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,111.5,-115,111.5</points>
<connection>
<GID>770</GID>
<name>IN_7</name></connection>
<connection>
<GID>786</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>24 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,107.5,-32,107.5</points>
<connection>
<GID>745</GID>
<name>IN_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>893 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,127.5,75,128.5</points>
<intersection>127.5 3</intersection>
<intersection>128.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,128.5,75,128.5</points>
<connection>
<GID>746</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75,127.5,75.5,127.5</points>
<connection>
<GID>743</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-128,55,-126.5,55</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<connection>
<GID>972</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1072 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,101.5,-25,101.5</points>
<connection>
<GID>761</GID>
<name>IN_0</name></connection>
<connection>
<GID>772</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1071 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-26,99.5,-25,99.5</points>
<connection>
<GID>761</GID>
<name>IN_1</name></connection>
<connection>
<GID>767</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1070 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18.5,100.5,-18.5,111</points>
<intersection>100.5 1</intersection>
<intersection>111 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-19,100.5,-18.5,100.5</points>
<connection>
<GID>761</GID>
<name>OUT</name></connection>
<intersection>-18.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-18.5,111,-18,111</points>
<connection>
<GID>549</GID>
<name>IN_2</name></connection>
<intersection>-18.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>918 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,103.5,-115,103.5</points>
<connection>
<GID>796</GID>
<name>IN_0</name></connection>
<connection>
<GID>774</GID>
<name>IN_7</name></connection></hsegment></shape></wire>
<wire>
<ID>919 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,107.5,-115,107.5</points>
<connection>
<GID>790</GID>
<name>IN_0</name></connection>
<connection>
<GID>774</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1094 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,47,135.5,47</points>
<connection>
<GID>765</GID>
<name>IN_0</name></connection>
<connection>
<GID>897</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1104 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,66,28,66</points>
<connection>
<GID>941</GID>
<name>IN_1</name></connection>
<connection>
<GID>943</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>925 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,52,21,52</points>
<connection>
<GID>794</GID>
<name>IN_0</name></connection>
<connection>
<GID>792</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>931 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,129,125.5,129</points>
<connection>
<GID>800</GID>
<name>IN_0</name></connection>
<connection>
<GID>802</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>992 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125,122.5,125,127</points>
<intersection>122.5 1</intersection>
<intersection>127 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,122.5,125,122.5</points>
<connection>
<GID>868</GID>
<name>OUT</name></connection>
<intersection>125 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125,127,125.5,127</points>
<connection>
<GID>800</GID>
<name>IN_1</name></connection>
<intersection>125 0</intersection></hsegment></shape></wire>
<wire>
<ID>1171 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,20.5,-75.5,20.5</points>
<connection>
<GID>1025</GID>
<name>IN_2</name></connection>
<connection>
<GID>1039</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>994 </ID>
<shape>
<hsegment>
<ID>13</ID>
<points>116.5,125.5,117.5,125.5</points>
<connection>
<GID>806</GID>
<name>IN_0</name></connection>
<connection>
<GID>868</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>993 </ID>
<shape>
<hsegment>
<ID>13</ID>
<points>116.5,123.5,117.5,123.5</points>
<connection>
<GID>808</GID>
<name>IN_0</name></connection>
<connection>
<GID>868</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>935 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19.5,39.5,21,39.5</points>
<connection>
<GID>810</GID>
<name>IN_0</name></connection>
<connection>
<GID>809</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1154 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-78,5.5,-78,8.5</points>
<intersection>5.5 2</intersection>
<intersection>8.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-78,8.5,-75.5,8.5</points>
<connection>
<GID>377</GID>
<name>IN_2</name></connection>
<intersection>-78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80,5.5,-78,5.5</points>
<connection>
<GID>775</GID>
<name>OUT</name></connection>
<intersection>-78 0</intersection></hsegment></shape></wire>
<wire>
<ID>947 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>91.5,5,92.5,5</points>
<connection>
<GID>817</GID>
<name>IN_0</name></connection>
<connection>
<GID>824</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1001 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,21,64,21</points>
<connection>
<GID>822</GID>
<name>IN_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1178 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,14.5,83.5,14.5</points>
<connection>
<GID>1050</GID>
<name>OUT</name></connection>
<intersection>83.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>83.5,7.5,83.5,14.5</points>
<intersection>7.5 5</intersection>
<intersection>14.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>83.5,7.5,84.5,7.5</points>
<connection>
<GID>824</GID>
<name>IN_1</name></connection>
<intersection>83.5 4</intersection></hsegment></shape></wire>
<wire>
<ID>1188 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>83,5.5,84.5,5.5</points>
<connection>
<GID>824</GID>
<name>IN_3</name></connection>
<connection>
<GID>1065</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1062 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-4.5,84,1.5</points>
<connection>
<GID>1072</GID>
<name>OUT_0</name></connection>
<intersection>1.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,1.5,84.5,1.5</points>
<connection>
<GID>824</GID>
<name>IN_4</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>1063 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>83.5,-4.5,83.5,2.5</points>
<intersection>-4.5 2</intersection>
<intersection>2.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,2.5,84.5,2.5</points>
<connection>
<GID>824</GID>
<name>IN_5</name></connection>
<intersection>83.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-4.5,83.5,-4.5</points>
<connection>
<GID>1073</GID>
<name>IN_0</name></connection>
<intersection>83.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1191 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82.5,1.5,82.5,4.5</points>
<intersection>1.5 2</intersection>
<intersection>4.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,4.5,84.5,4.5</points>
<connection>
<GID>824</GID>
<name>IN_7</name></connection>
<intersection>82.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,1.5,82.5,1.5</points>
<connection>
<GID>1069</GID>
<name>IN_0</name></connection>
<intersection>82.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1202 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,27.5,-86,27.5</points>
<connection>
<GID>1029</GID>
<name>IN_1</name></connection>
<connection>
<GID>1022</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1000 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>63,19,64,19</points>
<connection>
<GID>829</GID>
<name>IN_0</name></connection>
<connection>
<GID>875</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>960 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,118,-70,118</points>
<connection>
<GID>836</GID>
<name>IN_0</name></connection>
<connection>
<GID>838</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>961 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,116,-70,116</points>
<connection>
<GID>836</GID>
<name>IN_1</name></connection>
<connection>
<GID>840</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>943 </ID>
<shape>
<hsegment>
<ID>11</ID>
<points>-127.5,16,-126.5,16</points>
<connection>
<GID>845</GID>
<name>IN_0</name></connection>
<connection>
<GID>826</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>995 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,121.5,117.5,121.5</points>
<connection>
<GID>868</GID>
<name>IN_2</name></connection>
<connection>
<GID>869</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1145 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-133.5,2.5,-132.5,2.5</points>
<connection>
<GID>1008</GID>
<name>IN_0</name></connection>
<connection>
<GID>1002</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>996 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>116.5,119.5,117.5,119.5</points>
<connection>
<GID>868</GID>
<name>IN_3</name></connection>
<connection>
<GID>870</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>998 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,105,-70,105</points>
<connection>
<GID>871</GID>
<name>IN_1</name></connection>
<connection>
<GID>873</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,10,20,10</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<connection>
<GID>51</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1056 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,53.5,62,53.5</points>
<connection>
<GID>934</GID>
<name>IN_0</name></connection>
<connection>
<GID>937</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1055 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>61,51.5,62,51.5</points>
<connection>
<GID>934</GID>
<name>IN_1</name></connection>
<connection>
<GID>938</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1051 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>68,52.5,68,54</points>
<connection>
<GID>934</GID>
<name>OUT</name></connection>
<intersection>54 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68,54,68.5,54</points>
<connection>
<GID>931</GID>
<name>IN_1</name></connection>
<intersection>68 0</intersection></hsegment></shape></wire>
<wire>
<ID>1045 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>74.5,59.5,75.5,59.5</points>
<connection>
<GID>922</GID>
<name>IN_0</name></connection>
<connection>
<GID>904</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>18 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>12,4,13,4</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>19,2,20,2</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>1080 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,92,-19,92</points>
<connection>
<GID>881</GID>
<name>IN_0</name></connection>
<connection>
<GID>879</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1034 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>74.5,87.5,75.5,87.5</points>
<connection>
<GID>912</GID>
<name>IN_0</name></connection>
<connection>
<GID>899</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1083 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,83,-26,83</points>
<connection>
<GID>885</GID>
<name>IN_0</name></connection>
<connection>
<GID>884</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>86 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,19,130,19</points>
<connection>
<GID>618</GID>
<name>IN_0</name></connection>
<intersection>130 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130,19,130,19</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>19 1</intersection></vsegment></shape></wire>
<wire>
<ID>1082 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-27,81,-26,81</points>
<connection>
<GID>885</GID>
<name>IN_1</name></connection>
<connection>
<GID>883</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>81 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,-4,-126.5,-4</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>928 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,100.5,-115,100.5</points>
<connection>
<GID>799</GID>
<name>IN_0</name></connection>
<connection>
<GID>774</GID>
<name>IN_4</name></connection></hsegment></shape></wire>
<wire>
<ID>902 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,109.5,-32,109.5</points>
<connection>
<GID>733</GID>
<name>IN_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>27 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,100.5,-63,100.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71,101.5,-70,101.5</points>
<connection>
<GID>253</GID>
<name>IN_0</name></connection>
<connection>
<GID>255</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>946 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,96,121,96</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<connection>
<GID>300</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1123 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-135,56,-134,56</points>
<connection>
<GID>972</GID>
<name>IN_0</name></connection>
<connection>
<GID>971</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1124 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-135,54,-134,54</points>
<connection>
<GID>972</GID>
<name>IN_1</name></connection>
<connection>
<GID>973</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1142 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-69,16.5,-69,21.5</points>
<intersection>16.5 2</intersection>
<intersection>21.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-69,21.5,-68,21.5</points>
<connection>
<GID>755</GID>
<name>IN_1</name></connection>
<intersection>-69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,16.5,-69,16.5</points>
<connection>
<GID>757</GID>
<name>OUT</name></connection>
<intersection>-69 0</intersection></hsegment></shape></wire>
<wire>
<ID>321 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-71,94,-70,94</points>
<connection>
<GID>263</GID>
<name>IN_1</name></connection>
<connection>
<GID>265</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1119 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-127.5,41.5,-126.5,41.5</points>
<connection>
<GID>967</GID>
<name>IN_0</name></connection>
<connection>
<GID>965</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1169 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,24.5,-75.5,24.5</points>
<connection>
<GID>1025</GID>
<name>IN_0</name></connection>
<connection>
<GID>1037</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>326 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-64,89.5,-63,89.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<connection>
<GID>273</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>894 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>67.5,129.5,68.5,129.5</points>
<connection>
<GID>746</GID>
<name>IN_0</name></connection>
<connection>
<GID>747</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>895 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67.5,127.5,68.5,127.5</points>
<connection>
<GID>746</GID>
<name>IN_1</name></connection>
<connection>
<GID>749</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>323 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-71,90.5,-70,90.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<connection>
<GID>273</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1125 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,62,-126.5,62</points>
<connection>
<GID>975</GID>
<name>IN_0</name></connection>
<connection>
<GID>974</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1126 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,60,-126.5,60</points>
<connection>
<GID>975</GID>
<name>IN_1</name></connection>
<connection>
<GID>976</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1136 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-84,56.5,-83,56.5</points>
<connection>
<GID>980</GID>
<name>IN_1</name></connection>
<connection>
<GID>989</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>957 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>68,112,69,112</points>
<connection>
<GID>963</GID>
<name>IN_0</name></connection>
<connection>
<GID>960</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1140 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-126.5,3.5,-119.5,3.5</points>
<connection>
<GID>289</GID>
<name>J</name></connection>
<connection>
<GID>1002</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>83 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-120,-3,-120,-0.5</points>
<intersection>-3 2</intersection>
<intersection>-0.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-120,-0.5,-119.5,-0.5</points>
<connection>
<GID>289</GID>
<name>K</name></connection>
<intersection>-120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-120.5,-3,-120,-3</points>
<connection>
<GID>1</GID>
<name>OUT</name></connection>
<intersection>-120 0</intersection></hsegment></shape></wire>
<wire>
<ID>1110 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,67,21,67</points>
<connection>
<GID>943</GID>
<name>IN_0</name></connection>
<connection>
<GID>955</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>417 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,3.5,-111.5,3.5</points>
<connection>
<GID>289</GID>
<name>Q</name></connection>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>-112.5 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-112.5,3.5,-112.5,5</points>
<connection>
<GID>293</GID>
<name>N_in2</name></connection>
<intersection>3.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>955 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,106,27.5,108</points>
<intersection>106 1</intersection>
<intersection>108 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,106,27.5,106</points>
<connection>
<GID>548</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,108,28,108</points>
<connection>
<GID>930</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1162 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-92,-0.5,-91,-0.5</points>
<connection>
<GID>991</GID>
<name>IN_0</name></connection>
<connection>
<GID>992</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1172 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,-0.5,-86,-0.5</points>
<connection>
<GID>991</GID>
<name>OUT_0</name></connection>
<connection>
<GID>811</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>908 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-80,10.5,-75.5,10.5</points>
<connection>
<GID>671</GID>
<name>OUT</name></connection>
<connection>
<GID>377</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1057 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>134.5,90.5,135.5,90.5</points>
<connection>
<GID>979</GID>
<name>IN_0</name></connection>
<connection>
<GID>697</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>418 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,24,-53,24</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<connection>
<GID>297</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>1060 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-61.5,21.5,-61.5,24</points>
<intersection>21.5 2</intersection>
<intersection>24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-61.5,24,-61,24</points>
<connection>
<GID>297</GID>
<name>K</name></connection>
<intersection>-61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-62,21.5,-61.5,21.5</points>
<connection>
<GID>755</GID>
<name>OUT</name></connection>
<intersection>-61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>444 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-55,28,-53,28</points>
<connection>
<GID>297</GID>
<name>Q</name></connection>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-54 10</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>-54,28,-54,29.5</points>
<connection>
<GID>299</GID>
<name>N_in2</name></connection>
<intersection>28 1</intersection></vsegment></shape></wire>
<wire>
<ID>884 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,100,127.5,101</points>
<intersection>100 2</intersection>
<intersection>101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127,101,127.5,101</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,100,128,100</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>761 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,120,27.5,123</points>
<intersection>120 1</intersection>
<intersection>123 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,120,27.5,120</points>
<connection>
<GID>513</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,123,28,123</points>
<connection>
<GID>430</GID>
<name>IN_1</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>786 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>127.5,97,127.5,98</points>
<intersection>97 2</intersection>
<intersection>98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>127.5,98,128,98</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>127.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127,97,127.5,97</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>127.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1014 </ID>
<shape>
<hsegment>
<ID>17</ID>
<points>127.5,70,128.5,70</points>
<connection>
<GID>512</GID>
<name>IN_0</name></connection>
<connection>
<GID>485</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1144 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>-133.5,4.5,-132.5,4.5</points>
<connection>
<GID>1007</GID>
<name>IN_0</name></connection>
<connection>
<GID>1002</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1137 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11,13,-10,13</points>
<connection>
<GID>998</GID>
<name>IN_0</name></connection>
<connection>
<GID>995</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1116 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,46,-119.5,46</points>
<connection>
<GID>311</GID>
<name>J</name></connection>
<connection>
<GID>962</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>760 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,127.5,13.5,127.5</points>
<connection>
<GID>511</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-120,40.5,-120,42</points>
<intersection>40.5 2</intersection>
<intersection>42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-120,42,-119.5,42</points>
<connection>
<GID>311</GID>
<name>K</name></connection>
<intersection>-120 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-120.5,40.5,-120,40.5</points>
<connection>
<GID>965</GID>
<name>OUT</name></connection>
<intersection>-120 0</intersection></hsegment></shape></wire>
<wire>
<ID>1151 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-147.5,5.5,-146.5,5.5</points>
<connection>
<GID>1015</GID>
<name>IN_0</name></connection>
<connection>
<GID>1017</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1150 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-147.5,3.5,-146.5,3.5</points>
<connection>
<GID>1015</GID>
<name>IN_1</name></connection>
<connection>
<GID>1016</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-140,4.5,-140,7</points>
<intersection>4.5 1</intersection>
<intersection>7 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-140.5,4.5,-140,4.5</points>
<connection>
<GID>1015</GID>
<name>OUT</name></connection>
<intersection>-140 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-140,7,-139.5,7</points>
<connection>
<GID>1004</GID>
<name>IN_1</name></connection>
<intersection>-140 0</intersection></hsegment></shape></wire>
<wire>
<ID>709 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-113.5,29.5,-111.5,29.5</points>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<connection>
<GID>319</GID>
<name>nQ</name></connection></hsegment></shape></wire>
<wire>
<ID>1117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-120,28,-120,29.5</points>
<intersection>28 3</intersection>
<intersection>29.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-120,29.5,-119.5,29.5</points>
<connection>
<GID>319</GID>
<name>K</name></connection>
<intersection>-120 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-120.5,28,-120,28</points>
<connection>
<GID>964</GID>
<name>OUT</name></connection>
<intersection>-120 0</intersection></hsegment></shape></wire>
<wire>
<ID>1109 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,70,21,70</points>
<connection>
<GID>945</GID>
<name>IN_1</name></connection>
<connection>
<GID>954</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>759 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,129.5,13.5,129.5</points>
<connection>
<GID>484</GID>
<name>IN_0</name></connection>
<connection>
<GID>403</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1076 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,124.5,-32,124.5</points>
<connection>
<GID>814</GID>
<name>IN_0</name></connection>
<connection>
<GID>831</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1077 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,122.5,-32,122.5</points>
<connection>
<GID>814</GID>
<name>IN_1</name></connection>
<connection>
<GID>832</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1075 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,120.5,-32,120.5</points>
<connection>
<GID>814</GID>
<name>IN_2</name></connection>
<connection>
<GID>830</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>765 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,122,21,122</points>
<connection>
<GID>519</GID>
<name>IN_0</name></connection>
<connection>
<GID>513</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>766 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,120,21,120</points>
<connection>
<GID>521</GID>
<name>IN_0</name></connection>
<connection>
<GID>513</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>785 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,118,21,118</points>
<connection>
<GID>525</GID>
<name>IN_0</name></connection>
<connection>
<GID>513</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>1048 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,83.5,75.5,83.5</points>
<connection>
<GID>899</GID>
<name>IN_2</name></connection>
<connection>
<GID>927</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1122 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,27,-126.5,27</points>
<connection>
<GID>964</GID>
<name>IN_1</name></connection>
<connection>
<GID>970</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>787 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,107,21,107</points>
<connection>
<GID>552</GID>
<name>IN_0</name></connection>
<connection>
<GID>548</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1042 </ID>
<shape>
<hsegment>
<ID>5</ID>
<points>74.5,76.5,75.5,76.5</points>
<connection>
<GID>919</GID>
<name>IN_0</name></connection>
<connection>
<GID>900</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>881 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>27,99,28,99</points>
<connection>
<GID>595</GID>
<name>IN_1</name></connection>
<connection>
<GID>591</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>887 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,90.5,27.5,91.5</points>
<intersection>90.5 2</intersection>
<intersection>91.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,91.5,27.5,91.5</points>
<connection>
<GID>645</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,90.5,28,90.5</points>
<connection>
<GID>619</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>920 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,101.5,-115,101.5</points>
<connection>
<GID>798</GID>
<name>IN_0</name></connection>
<connection>
<GID>774</GID>
<name>IN_5</name></connection></hsegment></shape></wire>
<wire>
<ID>1093 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,46,128.5,46</points>
<connection>
<GID>897</GID>
<name>IN_1</name></connection>
<connection>
<GID>903</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>888 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>20,92.5,21,92.5</points>
<connection>
<GID>672</GID>
<name>IN_0</name></connection>
<connection>
<GID>645</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>889 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,90.5,21,90.5</points>
<connection>
<GID>676</GID>
<name>IN_0</name></connection>
<connection>
<GID>645</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1018 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,113,-18,113</points>
<connection>
<GID>623</GID>
<name>OUT</name></connection>
<connection>
<GID>549</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,34.5,-86,34.5</points>
<connection>
<GID>1030</GID>
<name>IN_0</name></connection>
<connection>
<GID>1028</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1027 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,104.5,75.5,104.5</points>
<connection>
<GID>894</GID>
<name>IN_0</name></connection>
<connection>
<GID>906</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1028 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,102.5,75.5,102.5</points>
<connection>
<GID>894</GID>
<name>IN_1</name></connection>
<connection>
<GID>905</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>897 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>67.5,123.5,68.5,123.5</points>
<connection>
<GID>741</GID>
<name>IN_1</name></connection>
<connection>
<GID>753</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>892 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,124.5,75,125.5</points>
<intersection>124.5 2</intersection>
<intersection>125.5 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>74.5,124.5,75,124.5</points>
<connection>
<GID>741</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75,125.5,75.5,125.5</points>
<connection>
<GID>743</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>1085 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,76,-19,76</points>
<connection>
<GID>888</GID>
<name>IN_1</name></connection>
<connection>
<GID>886</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>901 </ID>
<shape>
<hsegment>
<ID>23</ID>
<points>120,98,121,98</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1112 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,61.5,14,61.5</points>
<connection>
<GID>951</GID>
<name>IN_1</name></connection>
<connection>
<GID>957</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>933 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-124,104.5,-115,104.5</points>
<connection>
<GID>774</GID>
<name>IN_3</name></connection>
<connection>
<GID>795</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1061 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,22.5,-68.5,23.5</points>
<intersection>22.5 2</intersection>
<intersection>23.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,23.5,-68,23.5</points>
<connection>
<GID>755</GID>
<name>IN_0</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,22.5,-68.5,22.5</points>
<connection>
<GID>1025</GID>
<name>OUT</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-68.5,9.5,-68.5,19.5</points>
<intersection>9.5 2</intersection>
<intersection>19.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-68.5,19.5,-68,19.5</points>
<connection>
<GID>755</GID>
<name>IN_2</name></connection>
<intersection>-68.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-69.5,9.5,-68.5,9.5</points>
<connection>
<GID>377</GID>
<name>OUT</name></connection>
<intersection>-68.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1147 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,15.5,-75.5,15.5</points>
<connection>
<GID>757</GID>
<name>IN_1</name></connection>
<connection>
<GID>1044</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>944 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,90,-108,93</points>
<connection>
<GID>805</GID>
<name>OUT</name></connection>
<intersection>90 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,90,-107,90</points>
<connection>
<GID>804</GID>
<name>IN_0</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>945 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-108,85,-108,88</points>
<connection>
<GID>807</GID>
<name>OUT</name></connection>
<intersection>88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-108,88,-107,88</points>
<connection>
<GID>804</GID>
<name>IN_1</name></connection>
<intersection>-108 0</intersection></hsegment></shape></wire>
<wire>
<ID>1007 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-101,89,-100,89</points>
<connection>
<GID>804</GID>
<name>OUT</name></connection>
<connection>
<GID>878</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>965 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,96.5,-115,96.5</points>
<connection>
<GID>805</GID>
<name>IN_0</name></connection>
<connection>
<GID>816</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>983 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,95.5,-115,95.5</points>
<connection>
<GID>805</GID>
<name>IN_1</name></connection>
<connection>
<GID>818</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>982 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,93.5,-115,93.5</points>
<connection>
<GID>805</GID>
<name>IN_3</name></connection>
<connection>
<GID>825</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>977 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,90.5,-115,90.5</points>
<connection>
<GID>805</GID>
<name>IN_5</name></connection>
<connection>
<GID>835</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>976 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,92.5,-115,92.5</points>
<connection>
<GID>805</GID>
<name>IN_7</name></connection>
<connection>
<GID>827</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>951 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,88.5,-115,88.5</points>
<connection>
<GID>807</GID>
<name>IN_0</name></connection>
<connection>
<GID>839</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1157 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-77.5,0.5,-77.5,6.5</points>
<intersection>0.5 2</intersection>
<intersection>6.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-77.5,6.5,-75.5,6.5</points>
<connection>
<GID>377</GID>
<name>IN_3</name></connection>
<intersection>-77.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-80,0.5,-77.5,0.5</points>
<connection>
<GID>811</GID>
<name>OUT</name></connection>
<intersection>-77.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>952 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,86.5,-115,86.5</points>
<connection>
<GID>807</GID>
<name>IN_2</name></connection>
<connection>
<GID>846</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>979 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-125.5,81.5,-115,81.5</points>
<connection>
<GID>807</GID>
<name>IN_4</name></connection>
<connection>
<GID>874</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>953 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-116,82.5,-115,82.5</points>
<connection>
<GID>807</GID>
<name>IN_5</name></connection>
<connection>
<GID>867</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>82 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,-2,-126.5,-2</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<connection>
<GID>1</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1029 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,97.5,75.5,97.5</points>
<connection>
<GID>896</GID>
<name>IN_1</name></connection>
<connection>
<GID>907</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1031 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,94.5,75.5,94.5</points>
<connection>
<GID>898</GID>
<name>IN_0</name></connection>
<connection>
<GID>909</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1012 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,73.5,128.5,73.5</points>
<connection>
<GID>404</GID>
<name>IN_1</name></connection>
<connection>
<GID>458</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1033 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,92.5,75.5,92.5</points>
<connection>
<GID>898</GID>
<name>IN_1</name></connection>
<connection>
<GID>911</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1032 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,90.5,75.5,90.5</points>
<connection>
<GID>898</GID>
<name>IN_2</name></connection>
<connection>
<GID>910</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1038 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,73.5,75.5,73.5</points>
<connection>
<GID>901</GID>
<name>IN_0</name></connection>
<connection>
<GID>918</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1040 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,66.5,75.5,66.5</points>
<connection>
<GID>902</GID>
<name>IN_0</name></connection>
<connection>
<GID>920</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1047 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,64.5,75.5,64.5</points>
<connection>
<GID>902</GID>
<name>IN_1</name></connection>
<connection>
<GID>924</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1050 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,55,75,57.5</points>
<intersection>55 2</intersection>
<intersection>57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,57.5,75.5,57.5</points>
<connection>
<GID>904</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,55,75,55</points>
<connection>
<GID>931</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>1190 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,6.5,77,6.5</points>
<connection>
<GID>1065</GID>
<name>IN_0</name></connection>
<connection>
<GID>1066</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1066 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,43.5,69,43.5</points>
<connection>
<GID>944</GID>
<name>IN_0</name></connection>
<connection>
<GID>949</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1069 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,42.5,75,43.5</points>
<connection>
<GID>944</GID>
<name>OUT</name></connection>
<intersection>43.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>75,43.5,75.5,43.5</points>
<connection>
<GID>952</GID>
<name>IN_1</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>1068 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,45.5,75,46.5</points>
<intersection>45.5 3</intersection>
<intersection>46.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74,46.5,75,46.5</points>
<connection>
<GID>948</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75,45.5,75.5,45.5</points>
<connection>
<GID>952</GID>
<name>IN_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>413 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,111.5,128.5,111.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<connection>
<GID>56</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>681 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,109.5,128.5,109.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<connection>
<GID>60</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>899 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>120,100,121,100</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<connection>
<GID>285</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1011 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,75.5,128.5,75.5</points>
<connection>
<GID>404</GID>
<name>IN_0</name></connection>
<connection>
<GID>431</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>906 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,109.5,-25.5,112</points>
<intersection>109.5 2</intersection>
<intersection>112 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25.5,112,-25,112</points>
<connection>
<GID>623</GID>
<name>IN_1</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-26,109.5,-25.5,109.5</points>
<connection>
<GID>350</GID>
<name>OUT</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1015 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>127.5,68,128.5,68</points>
<connection>
<GID>485</GID>
<name>IN_1</name></connection>
<connection>
<GID>515</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1182 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,13.5,77,13.5</points>
<connection>
<GID>1054</GID>
<name>IN_0</name></connection>
<connection>
<GID>1050</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>905 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-33,111.5,-32,111.5</points>
<connection>
<GID>724</GID>
<name>IN_0</name></connection>
<connection>
<GID>350</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1106 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,68,27.5,71</points>
<intersection>68 1</intersection>
<intersection>71 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27.5,68,28,68</points>
<connection>
<GID>941</GID>
<name>IN_0</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27,71,27.5,71</points>
<connection>
<GID>945</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1105 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>27.5,57.5,27.5,64</points>
<intersection>57.5 1</intersection>
<intersection>64 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>27,57.5,27.5,57.5</points>
<connection>
<GID>946</GID>
<name>OUT</name></connection>
<intersection>27.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>27.5,64,28,64</points>
<connection>
<GID>941</GID>
<name>IN_2</name></connection>
<intersection>27.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1108 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,72,21,72</points>
<connection>
<GID>945</GID>
<name>IN_0</name></connection>
<connection>
<GID>953</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1114 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,56.5,21,56.5</points>
<connection>
<GID>959</GID>
<name>IN_0</name></connection>
<connection>
<GID>946</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>1111 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,63.5,14,63.5</points>
<connection>
<GID>951</GID>
<name>IN_0</name></connection>
<connection>
<GID>956</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1121 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,29,-126.5,29</points>
<connection>
<GID>964</GID>
<name>IN_0</name></connection>
<connection>
<GID>969</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1134 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-76.5,53,-76.5,60</points>
<intersection>53 3</intersection>
<intersection>57.5 2</intersection>
<intersection>60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-76.5,60,-73,60</points>
<connection>
<GID>982</GID>
<name>IN_1</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-77,57.5,-76.5,57.5</points>
<connection>
<GID>980</GID>
<name>OUT</name></connection>
<intersection>-76.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-76.5,53,-73,53</points>
<connection>
<GID>984</GID>
<name>IN_1</name></connection>
<intersection>-76.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-75,55,-75,55.5</points>
<connection>
<GID>986</GID>
<name>OUT_0</name></connection>
<intersection>55 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-75,55,-73,55</points>
<connection>
<GID>984</GID>
<name>IN_0</name></connection>
<intersection>-75 0</intersection></hsegment></shape></wire>
<wire>
<ID>1141 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-133,6.5,-133,8</points>
<intersection>6.5 2</intersection>
<intersection>8 3</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-133,6.5,-132.5,6.5</points>
<connection>
<GID>1002</GID>
<name>IN_0</name></connection>
<intersection>-133 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-133.5,8,-133,8</points>
<connection>
<GID>1004</GID>
<name>OUT</name></connection>
<intersection>-133 0</intersection></hsegment></shape></wire>
<wire>
<ID>1146 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>-133.5,0.5,-132.5,0.5</points>
<connection>
<GID>1002</GID>
<name>IN_3</name></connection>
<connection>
<GID>1009</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1152 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-140.5,9,-139.5,9</points>
<connection>
<GID>1004</GID>
<name>IN_0</name></connection>
<connection>
<GID>1018</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1170 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,22.5,-75.5,22.5</points>
<connection>
<GID>1025</GID>
<name>IN_1</name></connection>
<connection>
<GID>1038</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1164 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,46.5,-75.5,46.5</points>
<connection>
<GID>1023</GID>
<name>IN_1</name></connection>
<connection>
<GID>1032</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1165 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-76.5,44.5,-75.5,44.5</points>
<connection>
<GID>1023</GID>
<name>IN_2</name></connection>
<connection>
<GID>1033</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76,15.5,77,15.5</points>
<connection>
<GID>1050</GID>
<name>IN_0</name></connection>
<connection>
<GID>1052</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>937 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,20.5,-119.5,20.5</points>
<connection>
<GID>675</GID>
<name>J</name></connection>
<connection>
<GID>773</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>940 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-120,15,-120,16.5</points>
<intersection>15 3</intersection>
<intersection>16.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-120,16.5,-119.5,16.5</points>
<connection>
<GID>675</GID>
<name>K</name></connection>
<intersection>-120 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-120.5,15,-120,15</points>
<connection>
<GID>826</GID>
<name>OUT</name></connection>
<intersection>-120 0</intersection></hsegment></shape></wire>
<wire>
<ID>936 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-120.5,18.5,-119.5,18.5</points>
<connection>
<GID>675</GID>
<name>clock</name></connection>
<connection>
<GID>760</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>949 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-127.5,14,-126.5,14</points>
<connection>
<GID>826</GID>
<name>IN_1</name></connection>
<connection>
<GID>889</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>956 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,110,28,110</points>
<connection>
<GID>942</GID>
<name>IN_0</name></connection>
<connection>
<GID>930</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>958 </ID>
<shape>
<hsegment>
<ID>0</ID>
<points>68,110,69,110</points>
<connection>
<GID>947</GID>
<name>IN_0</name></connection>
<connection>
<GID>960</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>966 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,111,75.5,113</points>
<intersection>111 1</intersection>
<intersection>113 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,111,75.5,111</points>
<connection>
<GID>960</GID>
<name>OUT</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>75.5,113,76,113</points>
<connection>
<GID>966</GID>
<name>IN_1</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>1003 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,115,76,115</points>
<connection>
<GID>966</GID>
<name>IN_0</name></connection>
<connection>
<GID>977</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>1158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-87,6.5,-86,6.5</points>
<connection>
<GID>775</GID>
<name>IN_0</name></connection>
<connection>
<GID>834</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>87 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>129,17,130,17</points>
<connection>
<GID>754</GID>
<name>IN_0</name></connection>
<intersection>130 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>130,17,130,17</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>17 1</intersection></vsegment></shape></wire></page 2></circuit>